module RWSmem(
  input          clock,
  input          reset,
  input          io_enable,
  input          io_write,
  input  [6:0]   io_addr,
  input  [127:0] io_dataIn,
  output [127:0] io_dataOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [127:0] _RAND_27;
  reg [127:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [127:0] _RAND_33;
  reg [127:0] _RAND_34;
  reg [127:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [127:0] _RAND_38;
  reg [127:0] _RAND_39;
  reg [127:0] _RAND_40;
  reg [127:0] _RAND_41;
  reg [127:0] _RAND_42;
  reg [127:0] _RAND_43;
  reg [127:0] _RAND_44;
  reg [127:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [127:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [127:0] _RAND_50;
  reg [127:0] _RAND_51;
  reg [127:0] _RAND_52;
  reg [127:0] _RAND_53;
  reg [127:0] _RAND_54;
  reg [127:0] _RAND_55;
  reg [127:0] _RAND_56;
  reg [127:0] _RAND_57;
  reg [127:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [127:0] _RAND_61;
  reg [127:0] _RAND_62;
  reg [127:0] _RAND_63;
  reg [127:0] _RAND_64;
  reg [127:0] _RAND_65;
  reg [127:0] _RAND_66;
  reg [127:0] _RAND_67;
  reg [127:0] _RAND_68;
  reg [127:0] _RAND_69;
  reg [127:0] _RAND_70;
  reg [127:0] _RAND_71;
  reg [127:0] _RAND_72;
  reg [127:0] _RAND_73;
  reg [127:0] _RAND_74;
  reg [127:0] _RAND_75;
  reg [127:0] _RAND_76;
  reg [127:0] _RAND_77;
  reg [127:0] _RAND_78;
  reg [127:0] _RAND_79;
  reg [127:0] _RAND_80;
  reg [127:0] _RAND_81;
  reg [127:0] _RAND_82;
  reg [127:0] _RAND_83;
  reg [127:0] _RAND_84;
  reg [127:0] _RAND_85;
  reg [127:0] _RAND_86;
  reg [127:0] _RAND_87;
  reg [127:0] _RAND_88;
  reg [127:0] _RAND_89;
  reg [127:0] _RAND_90;
  reg [127:0] _RAND_91;
  reg [127:0] _RAND_92;
  reg [127:0] _RAND_93;
  reg [127:0] _RAND_94;
  reg [127:0] _RAND_95;
  reg [127:0] _RAND_96;
  reg [127:0] _RAND_97;
  reg [127:0] _RAND_98;
  reg [127:0] _RAND_99;
  reg [127:0] _RAND_100;
  reg [127:0] _RAND_101;
  reg [127:0] _RAND_102;
  reg [127:0] _RAND_103;
  reg [127:0] _RAND_104;
  reg [127:0] _RAND_105;
  reg [127:0] _RAND_106;
  reg [127:0] _RAND_107;
  reg [127:0] _RAND_108;
  reg [127:0] _RAND_109;
  reg [127:0] _RAND_110;
  reg [127:0] _RAND_111;
  reg [127:0] _RAND_112;
  reg [127:0] _RAND_113;
  reg [127:0] _RAND_114;
  reg [127:0] _RAND_115;
  reg [127:0] _RAND_116;
  reg [127:0] _RAND_117;
  reg [127:0] _RAND_118;
  reg [127:0] _RAND_119;
  reg [127:0] _RAND_120;
  reg [127:0] _RAND_121;
  reg [127:0] _RAND_122;
  reg [127:0] _RAND_123;
  reg [127:0] _RAND_124;
  reg [127:0] _RAND_125;
  reg [127:0] _RAND_126;
  reg [127:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] mem_0; // @[Ram.scala 16:16]
  reg [127:0] mem_1; // @[Ram.scala 16:16]
  reg [127:0] mem_2; // @[Ram.scala 16:16]
  reg [127:0] mem_3; // @[Ram.scala 16:16]
  reg [127:0] mem_4; // @[Ram.scala 16:16]
  reg [127:0] mem_5; // @[Ram.scala 16:16]
  reg [127:0] mem_6; // @[Ram.scala 16:16]
  reg [127:0] mem_7; // @[Ram.scala 16:16]
  reg [127:0] mem_8; // @[Ram.scala 16:16]
  reg [127:0] mem_9; // @[Ram.scala 16:16]
  reg [127:0] mem_10; // @[Ram.scala 16:16]
  reg [127:0] mem_11; // @[Ram.scala 16:16]
  reg [127:0] mem_12; // @[Ram.scala 16:16]
  reg [127:0] mem_13; // @[Ram.scala 16:16]
  reg [127:0] mem_14; // @[Ram.scala 16:16]
  reg [127:0] mem_15; // @[Ram.scala 16:16]
  reg [127:0] mem_16; // @[Ram.scala 16:16]
  reg [127:0] mem_17; // @[Ram.scala 16:16]
  reg [127:0] mem_18; // @[Ram.scala 16:16]
  reg [127:0] mem_19; // @[Ram.scala 16:16]
  reg [127:0] mem_20; // @[Ram.scala 16:16]
  reg [127:0] mem_21; // @[Ram.scala 16:16]
  reg [127:0] mem_22; // @[Ram.scala 16:16]
  reg [127:0] mem_23; // @[Ram.scala 16:16]
  reg [127:0] mem_24; // @[Ram.scala 16:16]
  reg [127:0] mem_25; // @[Ram.scala 16:16]
  reg [127:0] mem_26; // @[Ram.scala 16:16]
  reg [127:0] mem_27; // @[Ram.scala 16:16]
  reg [127:0] mem_28; // @[Ram.scala 16:16]
  reg [127:0] mem_29; // @[Ram.scala 16:16]
  reg [127:0] mem_30; // @[Ram.scala 16:16]
  reg [127:0] mem_31; // @[Ram.scala 16:16]
  reg [127:0] mem_32; // @[Ram.scala 16:16]
  reg [127:0] mem_33; // @[Ram.scala 16:16]
  reg [127:0] mem_34; // @[Ram.scala 16:16]
  reg [127:0] mem_35; // @[Ram.scala 16:16]
  reg [127:0] mem_36; // @[Ram.scala 16:16]
  reg [127:0] mem_37; // @[Ram.scala 16:16]
  reg [127:0] mem_38; // @[Ram.scala 16:16]
  reg [127:0] mem_39; // @[Ram.scala 16:16]
  reg [127:0] mem_40; // @[Ram.scala 16:16]
  reg [127:0] mem_41; // @[Ram.scala 16:16]
  reg [127:0] mem_42; // @[Ram.scala 16:16]
  reg [127:0] mem_43; // @[Ram.scala 16:16]
  reg [127:0] mem_44; // @[Ram.scala 16:16]
  reg [127:0] mem_45; // @[Ram.scala 16:16]
  reg [127:0] mem_46; // @[Ram.scala 16:16]
  reg [127:0] mem_47; // @[Ram.scala 16:16]
  reg [127:0] mem_48; // @[Ram.scala 16:16]
  reg [127:0] mem_49; // @[Ram.scala 16:16]
  reg [127:0] mem_50; // @[Ram.scala 16:16]
  reg [127:0] mem_51; // @[Ram.scala 16:16]
  reg [127:0] mem_52; // @[Ram.scala 16:16]
  reg [127:0] mem_53; // @[Ram.scala 16:16]
  reg [127:0] mem_54; // @[Ram.scala 16:16]
  reg [127:0] mem_55; // @[Ram.scala 16:16]
  reg [127:0] mem_56; // @[Ram.scala 16:16]
  reg [127:0] mem_57; // @[Ram.scala 16:16]
  reg [127:0] mem_58; // @[Ram.scala 16:16]
  reg [127:0] mem_59; // @[Ram.scala 16:16]
  reg [127:0] mem_60; // @[Ram.scala 16:16]
  reg [127:0] mem_61; // @[Ram.scala 16:16]
  reg [127:0] mem_62; // @[Ram.scala 16:16]
  reg [127:0] mem_63; // @[Ram.scala 16:16]
  reg [127:0] mem_64; // @[Ram.scala 16:16]
  reg [127:0] mem_65; // @[Ram.scala 16:16]
  reg [127:0] mem_66; // @[Ram.scala 16:16]
  reg [127:0] mem_67; // @[Ram.scala 16:16]
  reg [127:0] mem_68; // @[Ram.scala 16:16]
  reg [127:0] mem_69; // @[Ram.scala 16:16]
  reg [127:0] mem_70; // @[Ram.scala 16:16]
  reg [127:0] mem_71; // @[Ram.scala 16:16]
  reg [127:0] mem_72; // @[Ram.scala 16:16]
  reg [127:0] mem_73; // @[Ram.scala 16:16]
  reg [127:0] mem_74; // @[Ram.scala 16:16]
  reg [127:0] mem_75; // @[Ram.scala 16:16]
  reg [127:0] mem_76; // @[Ram.scala 16:16]
  reg [127:0] mem_77; // @[Ram.scala 16:16]
  reg [127:0] mem_78; // @[Ram.scala 16:16]
  reg [127:0] mem_79; // @[Ram.scala 16:16]
  reg [127:0] mem_80; // @[Ram.scala 16:16]
  reg [127:0] mem_81; // @[Ram.scala 16:16]
  reg [127:0] mem_82; // @[Ram.scala 16:16]
  reg [127:0] mem_83; // @[Ram.scala 16:16]
  reg [127:0] mem_84; // @[Ram.scala 16:16]
  reg [127:0] mem_85; // @[Ram.scala 16:16]
  reg [127:0] mem_86; // @[Ram.scala 16:16]
  reg [127:0] mem_87; // @[Ram.scala 16:16]
  reg [127:0] mem_88; // @[Ram.scala 16:16]
  reg [127:0] mem_89; // @[Ram.scala 16:16]
  reg [127:0] mem_90; // @[Ram.scala 16:16]
  reg [127:0] mem_91; // @[Ram.scala 16:16]
  reg [127:0] mem_92; // @[Ram.scala 16:16]
  reg [127:0] mem_93; // @[Ram.scala 16:16]
  reg [127:0] mem_94; // @[Ram.scala 16:16]
  reg [127:0] mem_95; // @[Ram.scala 16:16]
  reg [127:0] mem_96; // @[Ram.scala 16:16]
  reg [127:0] mem_97; // @[Ram.scala 16:16]
  reg [127:0] mem_98; // @[Ram.scala 16:16]
  reg [127:0] mem_99; // @[Ram.scala 16:16]
  reg [127:0] mem_100; // @[Ram.scala 16:16]
  reg [127:0] mem_101; // @[Ram.scala 16:16]
  reg [127:0] mem_102; // @[Ram.scala 16:16]
  reg [127:0] mem_103; // @[Ram.scala 16:16]
  reg [127:0] mem_104; // @[Ram.scala 16:16]
  reg [127:0] mem_105; // @[Ram.scala 16:16]
  reg [127:0] mem_106; // @[Ram.scala 16:16]
  reg [127:0] mem_107; // @[Ram.scala 16:16]
  reg [127:0] mem_108; // @[Ram.scala 16:16]
  reg [127:0] mem_109; // @[Ram.scala 16:16]
  reg [127:0] mem_110; // @[Ram.scala 16:16]
  reg [127:0] mem_111; // @[Ram.scala 16:16]
  reg [127:0] mem_112; // @[Ram.scala 16:16]
  reg [127:0] mem_113; // @[Ram.scala 16:16]
  reg [127:0] mem_114; // @[Ram.scala 16:16]
  reg [127:0] mem_115; // @[Ram.scala 16:16]
  reg [127:0] mem_116; // @[Ram.scala 16:16]
  reg [127:0] mem_117; // @[Ram.scala 16:16]
  reg [127:0] mem_118; // @[Ram.scala 16:16]
  reg [127:0] mem_119; // @[Ram.scala 16:16]
  reg [127:0] mem_120; // @[Ram.scala 16:16]
  reg [127:0] mem_121; // @[Ram.scala 16:16]
  reg [127:0] mem_122; // @[Ram.scala 16:16]
  reg [127:0] mem_123; // @[Ram.scala 16:16]
  reg [127:0] mem_124; // @[Ram.scala 16:16]
  reg [127:0] mem_125; // @[Ram.scala 16:16]
  reg [127:0] mem_126; // @[Ram.scala 16:16]
  reg [127:0] mem_127; // @[Ram.scala 16:16]
  wire [127:0] _GEN_129 = 7'h1 == io_addr ? mem_1 : mem_0; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_130 = 7'h2 == io_addr ? mem_2 : _GEN_129; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_131 = 7'h3 == io_addr ? mem_3 : _GEN_130; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_132 = 7'h4 == io_addr ? mem_4 : _GEN_131; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_133 = 7'h5 == io_addr ? mem_5 : _GEN_132; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_134 = 7'h6 == io_addr ? mem_6 : _GEN_133; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_135 = 7'h7 == io_addr ? mem_7 : _GEN_134; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_136 = 7'h8 == io_addr ? mem_8 : _GEN_135; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_137 = 7'h9 == io_addr ? mem_9 : _GEN_136; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_138 = 7'ha == io_addr ? mem_10 : _GEN_137; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_139 = 7'hb == io_addr ? mem_11 : _GEN_138; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_140 = 7'hc == io_addr ? mem_12 : _GEN_139; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_141 = 7'hd == io_addr ? mem_13 : _GEN_140; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_142 = 7'he == io_addr ? mem_14 : _GEN_141; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_143 = 7'hf == io_addr ? mem_15 : _GEN_142; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_144 = 7'h10 == io_addr ? mem_16 : _GEN_143; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_145 = 7'h11 == io_addr ? mem_17 : _GEN_144; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_146 = 7'h12 == io_addr ? mem_18 : _GEN_145; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_147 = 7'h13 == io_addr ? mem_19 : _GEN_146; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_148 = 7'h14 == io_addr ? mem_20 : _GEN_147; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_149 = 7'h15 == io_addr ? mem_21 : _GEN_148; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_150 = 7'h16 == io_addr ? mem_22 : _GEN_149; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_151 = 7'h17 == io_addr ? mem_23 : _GEN_150; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_152 = 7'h18 == io_addr ? mem_24 : _GEN_151; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_153 = 7'h19 == io_addr ? mem_25 : _GEN_152; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_154 = 7'h1a == io_addr ? mem_26 : _GEN_153; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_155 = 7'h1b == io_addr ? mem_27 : _GEN_154; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_156 = 7'h1c == io_addr ? mem_28 : _GEN_155; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_157 = 7'h1d == io_addr ? mem_29 : _GEN_156; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_158 = 7'h1e == io_addr ? mem_30 : _GEN_157; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_159 = 7'h1f == io_addr ? mem_31 : _GEN_158; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_160 = 7'h20 == io_addr ? mem_32 : _GEN_159; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_161 = 7'h21 == io_addr ? mem_33 : _GEN_160; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_162 = 7'h22 == io_addr ? mem_34 : _GEN_161; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_163 = 7'h23 == io_addr ? mem_35 : _GEN_162; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_164 = 7'h24 == io_addr ? mem_36 : _GEN_163; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_165 = 7'h25 == io_addr ? mem_37 : _GEN_164; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_166 = 7'h26 == io_addr ? mem_38 : _GEN_165; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_167 = 7'h27 == io_addr ? mem_39 : _GEN_166; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_168 = 7'h28 == io_addr ? mem_40 : _GEN_167; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_169 = 7'h29 == io_addr ? mem_41 : _GEN_168; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_170 = 7'h2a == io_addr ? mem_42 : _GEN_169; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_171 = 7'h2b == io_addr ? mem_43 : _GEN_170; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_172 = 7'h2c == io_addr ? mem_44 : _GEN_171; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_173 = 7'h2d == io_addr ? mem_45 : _GEN_172; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_174 = 7'h2e == io_addr ? mem_46 : _GEN_173; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_175 = 7'h2f == io_addr ? mem_47 : _GEN_174; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_176 = 7'h30 == io_addr ? mem_48 : _GEN_175; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_177 = 7'h31 == io_addr ? mem_49 : _GEN_176; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_178 = 7'h32 == io_addr ? mem_50 : _GEN_177; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_179 = 7'h33 == io_addr ? mem_51 : _GEN_178; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_180 = 7'h34 == io_addr ? mem_52 : _GEN_179; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_181 = 7'h35 == io_addr ? mem_53 : _GEN_180; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_182 = 7'h36 == io_addr ? mem_54 : _GEN_181; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_183 = 7'h37 == io_addr ? mem_55 : _GEN_182; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_184 = 7'h38 == io_addr ? mem_56 : _GEN_183; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_185 = 7'h39 == io_addr ? mem_57 : _GEN_184; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_186 = 7'h3a == io_addr ? mem_58 : _GEN_185; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_187 = 7'h3b == io_addr ? mem_59 : _GEN_186; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_188 = 7'h3c == io_addr ? mem_60 : _GEN_187; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_189 = 7'h3d == io_addr ? mem_61 : _GEN_188; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_190 = 7'h3e == io_addr ? mem_62 : _GEN_189; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_191 = 7'h3f == io_addr ? mem_63 : _GEN_190; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_192 = 7'h40 == io_addr ? mem_64 : _GEN_191; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_193 = 7'h41 == io_addr ? mem_65 : _GEN_192; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_194 = 7'h42 == io_addr ? mem_66 : _GEN_193; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_195 = 7'h43 == io_addr ? mem_67 : _GEN_194; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_196 = 7'h44 == io_addr ? mem_68 : _GEN_195; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_197 = 7'h45 == io_addr ? mem_69 : _GEN_196; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_198 = 7'h46 == io_addr ? mem_70 : _GEN_197; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_199 = 7'h47 == io_addr ? mem_71 : _GEN_198; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_200 = 7'h48 == io_addr ? mem_72 : _GEN_199; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_201 = 7'h49 == io_addr ? mem_73 : _GEN_200; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_202 = 7'h4a == io_addr ? mem_74 : _GEN_201; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_203 = 7'h4b == io_addr ? mem_75 : _GEN_202; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_204 = 7'h4c == io_addr ? mem_76 : _GEN_203; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_205 = 7'h4d == io_addr ? mem_77 : _GEN_204; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_206 = 7'h4e == io_addr ? mem_78 : _GEN_205; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_207 = 7'h4f == io_addr ? mem_79 : _GEN_206; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_208 = 7'h50 == io_addr ? mem_80 : _GEN_207; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_209 = 7'h51 == io_addr ? mem_81 : _GEN_208; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_210 = 7'h52 == io_addr ? mem_82 : _GEN_209; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_211 = 7'h53 == io_addr ? mem_83 : _GEN_210; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_212 = 7'h54 == io_addr ? mem_84 : _GEN_211; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_213 = 7'h55 == io_addr ? mem_85 : _GEN_212; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_214 = 7'h56 == io_addr ? mem_86 : _GEN_213; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_215 = 7'h57 == io_addr ? mem_87 : _GEN_214; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_216 = 7'h58 == io_addr ? mem_88 : _GEN_215; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_217 = 7'h59 == io_addr ? mem_89 : _GEN_216; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_218 = 7'h5a == io_addr ? mem_90 : _GEN_217; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_219 = 7'h5b == io_addr ? mem_91 : _GEN_218; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_220 = 7'h5c == io_addr ? mem_92 : _GEN_219; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_221 = 7'h5d == io_addr ? mem_93 : _GEN_220; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_222 = 7'h5e == io_addr ? mem_94 : _GEN_221; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_223 = 7'h5f == io_addr ? mem_95 : _GEN_222; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_224 = 7'h60 == io_addr ? mem_96 : _GEN_223; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_225 = 7'h61 == io_addr ? mem_97 : _GEN_224; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_226 = 7'h62 == io_addr ? mem_98 : _GEN_225; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_227 = 7'h63 == io_addr ? mem_99 : _GEN_226; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_228 = 7'h64 == io_addr ? mem_100 : _GEN_227; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_229 = 7'h65 == io_addr ? mem_101 : _GEN_228; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_230 = 7'h66 == io_addr ? mem_102 : _GEN_229; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_231 = 7'h67 == io_addr ? mem_103 : _GEN_230; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_232 = 7'h68 == io_addr ? mem_104 : _GEN_231; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_233 = 7'h69 == io_addr ? mem_105 : _GEN_232; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_234 = 7'h6a == io_addr ? mem_106 : _GEN_233; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_235 = 7'h6b == io_addr ? mem_107 : _GEN_234; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_236 = 7'h6c == io_addr ? mem_108 : _GEN_235; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_237 = 7'h6d == io_addr ? mem_109 : _GEN_236; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_238 = 7'h6e == io_addr ? mem_110 : _GEN_237; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_239 = 7'h6f == io_addr ? mem_111 : _GEN_238; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_240 = 7'h70 == io_addr ? mem_112 : _GEN_239; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_241 = 7'h71 == io_addr ? mem_113 : _GEN_240; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_242 = 7'h72 == io_addr ? mem_114 : _GEN_241; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_243 = 7'h73 == io_addr ? mem_115 : _GEN_242; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_244 = 7'h74 == io_addr ? mem_116 : _GEN_243; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_245 = 7'h75 == io_addr ? mem_117 : _GEN_244; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_246 = 7'h76 == io_addr ? mem_118 : _GEN_245; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_247 = 7'h77 == io_addr ? mem_119 : _GEN_246; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_248 = 7'h78 == io_addr ? mem_120 : _GEN_247; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_249 = 7'h79 == io_addr ? mem_121 : _GEN_248; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_250 = 7'h7a == io_addr ? mem_122 : _GEN_249; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_251 = 7'h7b == io_addr ? mem_123 : _GEN_250; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_252 = 7'h7c == io_addr ? mem_124 : _GEN_251; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_253 = 7'h7d == io_addr ? mem_125 : _GEN_252; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_254 = 7'h7e == io_addr ? mem_126 : _GEN_253; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_255 = 7'h7f == io_addr ? mem_127 : _GEN_254; // @[Ram.scala 20:{31,31}]
  wire [127:0] _GEN_384 = io_write ? 128'h0 : _GEN_255; // @[Ram.scala 17:14 19:20 20:31]
  assign io_dataOut = io_enable ? _GEN_384 : 128'h0; // @[Ram.scala 17:14 18:19]
  always @(posedge clock) begin
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h0 == io_addr) begin // @[Ram.scala 19:35]
          mem_0 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h1 == io_addr) begin // @[Ram.scala 19:35]
          mem_1 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h2 == io_addr) begin // @[Ram.scala 19:35]
          mem_2 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h3 == io_addr) begin // @[Ram.scala 19:35]
          mem_3 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h4 == io_addr) begin // @[Ram.scala 19:35]
          mem_4 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h5 == io_addr) begin // @[Ram.scala 19:35]
          mem_5 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h6 == io_addr) begin // @[Ram.scala 19:35]
          mem_6 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h7 == io_addr) begin // @[Ram.scala 19:35]
          mem_7 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h8 == io_addr) begin // @[Ram.scala 19:35]
          mem_8 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h9 == io_addr) begin // @[Ram.scala 19:35]
          mem_9 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'ha == io_addr) begin // @[Ram.scala 19:35]
          mem_10 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'hb == io_addr) begin // @[Ram.scala 19:35]
          mem_11 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'hc == io_addr) begin // @[Ram.scala 19:35]
          mem_12 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'hd == io_addr) begin // @[Ram.scala 19:35]
          mem_13 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'he == io_addr) begin // @[Ram.scala 19:35]
          mem_14 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'hf == io_addr) begin // @[Ram.scala 19:35]
          mem_15 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h10 == io_addr) begin // @[Ram.scala 19:35]
          mem_16 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h11 == io_addr) begin // @[Ram.scala 19:35]
          mem_17 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h12 == io_addr) begin // @[Ram.scala 19:35]
          mem_18 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h13 == io_addr) begin // @[Ram.scala 19:35]
          mem_19 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h14 == io_addr) begin // @[Ram.scala 19:35]
          mem_20 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h15 == io_addr) begin // @[Ram.scala 19:35]
          mem_21 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h16 == io_addr) begin // @[Ram.scala 19:35]
          mem_22 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h17 == io_addr) begin // @[Ram.scala 19:35]
          mem_23 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h18 == io_addr) begin // @[Ram.scala 19:35]
          mem_24 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h19 == io_addr) begin // @[Ram.scala 19:35]
          mem_25 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h1a == io_addr) begin // @[Ram.scala 19:35]
          mem_26 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h1b == io_addr) begin // @[Ram.scala 19:35]
          mem_27 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h1c == io_addr) begin // @[Ram.scala 19:35]
          mem_28 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h1d == io_addr) begin // @[Ram.scala 19:35]
          mem_29 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h1e == io_addr) begin // @[Ram.scala 19:35]
          mem_30 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h1f == io_addr) begin // @[Ram.scala 19:35]
          mem_31 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h20 == io_addr) begin // @[Ram.scala 19:35]
          mem_32 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h21 == io_addr) begin // @[Ram.scala 19:35]
          mem_33 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h22 == io_addr) begin // @[Ram.scala 19:35]
          mem_34 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h23 == io_addr) begin // @[Ram.scala 19:35]
          mem_35 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h24 == io_addr) begin // @[Ram.scala 19:35]
          mem_36 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h25 == io_addr) begin // @[Ram.scala 19:35]
          mem_37 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h26 == io_addr) begin // @[Ram.scala 19:35]
          mem_38 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h27 == io_addr) begin // @[Ram.scala 19:35]
          mem_39 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h28 == io_addr) begin // @[Ram.scala 19:35]
          mem_40 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h29 == io_addr) begin // @[Ram.scala 19:35]
          mem_41 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h2a == io_addr) begin // @[Ram.scala 19:35]
          mem_42 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h2b == io_addr) begin // @[Ram.scala 19:35]
          mem_43 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h2c == io_addr) begin // @[Ram.scala 19:35]
          mem_44 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h2d == io_addr) begin // @[Ram.scala 19:35]
          mem_45 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h2e == io_addr) begin // @[Ram.scala 19:35]
          mem_46 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h2f == io_addr) begin // @[Ram.scala 19:35]
          mem_47 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h30 == io_addr) begin // @[Ram.scala 19:35]
          mem_48 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h31 == io_addr) begin // @[Ram.scala 19:35]
          mem_49 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h32 == io_addr) begin // @[Ram.scala 19:35]
          mem_50 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h33 == io_addr) begin // @[Ram.scala 19:35]
          mem_51 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h34 == io_addr) begin // @[Ram.scala 19:35]
          mem_52 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h35 == io_addr) begin // @[Ram.scala 19:35]
          mem_53 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h36 == io_addr) begin // @[Ram.scala 19:35]
          mem_54 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h37 == io_addr) begin // @[Ram.scala 19:35]
          mem_55 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h38 == io_addr) begin // @[Ram.scala 19:35]
          mem_56 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h39 == io_addr) begin // @[Ram.scala 19:35]
          mem_57 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h3a == io_addr) begin // @[Ram.scala 19:35]
          mem_58 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h3b == io_addr) begin // @[Ram.scala 19:35]
          mem_59 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h3c == io_addr) begin // @[Ram.scala 19:35]
          mem_60 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h3d == io_addr) begin // @[Ram.scala 19:35]
          mem_61 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h3e == io_addr) begin // @[Ram.scala 19:35]
          mem_62 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h3f == io_addr) begin // @[Ram.scala 19:35]
          mem_63 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h40 == io_addr) begin // @[Ram.scala 19:35]
          mem_64 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h41 == io_addr) begin // @[Ram.scala 19:35]
          mem_65 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h42 == io_addr) begin // @[Ram.scala 19:35]
          mem_66 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h43 == io_addr) begin // @[Ram.scala 19:35]
          mem_67 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h44 == io_addr) begin // @[Ram.scala 19:35]
          mem_68 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h45 == io_addr) begin // @[Ram.scala 19:35]
          mem_69 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h46 == io_addr) begin // @[Ram.scala 19:35]
          mem_70 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h47 == io_addr) begin // @[Ram.scala 19:35]
          mem_71 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h48 == io_addr) begin // @[Ram.scala 19:35]
          mem_72 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h49 == io_addr) begin // @[Ram.scala 19:35]
          mem_73 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h4a == io_addr) begin // @[Ram.scala 19:35]
          mem_74 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h4b == io_addr) begin // @[Ram.scala 19:35]
          mem_75 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h4c == io_addr) begin // @[Ram.scala 19:35]
          mem_76 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h4d == io_addr) begin // @[Ram.scala 19:35]
          mem_77 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h4e == io_addr) begin // @[Ram.scala 19:35]
          mem_78 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h4f == io_addr) begin // @[Ram.scala 19:35]
          mem_79 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h50 == io_addr) begin // @[Ram.scala 19:35]
          mem_80 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h51 == io_addr) begin // @[Ram.scala 19:35]
          mem_81 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h52 == io_addr) begin // @[Ram.scala 19:35]
          mem_82 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h53 == io_addr) begin // @[Ram.scala 19:35]
          mem_83 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h54 == io_addr) begin // @[Ram.scala 19:35]
          mem_84 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h55 == io_addr) begin // @[Ram.scala 19:35]
          mem_85 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h56 == io_addr) begin // @[Ram.scala 19:35]
          mem_86 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h57 == io_addr) begin // @[Ram.scala 19:35]
          mem_87 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h58 == io_addr) begin // @[Ram.scala 19:35]
          mem_88 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h59 == io_addr) begin // @[Ram.scala 19:35]
          mem_89 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h5a == io_addr) begin // @[Ram.scala 19:35]
          mem_90 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h5b == io_addr) begin // @[Ram.scala 19:35]
          mem_91 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h5c == io_addr) begin // @[Ram.scala 19:35]
          mem_92 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h5d == io_addr) begin // @[Ram.scala 19:35]
          mem_93 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h5e == io_addr) begin // @[Ram.scala 19:35]
          mem_94 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h5f == io_addr) begin // @[Ram.scala 19:35]
          mem_95 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h60 == io_addr) begin // @[Ram.scala 19:35]
          mem_96 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h61 == io_addr) begin // @[Ram.scala 19:35]
          mem_97 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h62 == io_addr) begin // @[Ram.scala 19:35]
          mem_98 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h63 == io_addr) begin // @[Ram.scala 19:35]
          mem_99 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h64 == io_addr) begin // @[Ram.scala 19:35]
          mem_100 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h65 == io_addr) begin // @[Ram.scala 19:35]
          mem_101 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h66 == io_addr) begin // @[Ram.scala 19:35]
          mem_102 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h67 == io_addr) begin // @[Ram.scala 19:35]
          mem_103 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h68 == io_addr) begin // @[Ram.scala 19:35]
          mem_104 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h69 == io_addr) begin // @[Ram.scala 19:35]
          mem_105 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h6a == io_addr) begin // @[Ram.scala 19:35]
          mem_106 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h6b == io_addr) begin // @[Ram.scala 19:35]
          mem_107 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h6c == io_addr) begin // @[Ram.scala 19:35]
          mem_108 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h6d == io_addr) begin // @[Ram.scala 19:35]
          mem_109 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h6e == io_addr) begin // @[Ram.scala 19:35]
          mem_110 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h6f == io_addr) begin // @[Ram.scala 19:35]
          mem_111 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h70 == io_addr) begin // @[Ram.scala 19:35]
          mem_112 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h71 == io_addr) begin // @[Ram.scala 19:35]
          mem_113 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h72 == io_addr) begin // @[Ram.scala 19:35]
          mem_114 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h73 == io_addr) begin // @[Ram.scala 19:35]
          mem_115 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h74 == io_addr) begin // @[Ram.scala 19:35]
          mem_116 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h75 == io_addr) begin // @[Ram.scala 19:35]
          mem_117 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h76 == io_addr) begin // @[Ram.scala 19:35]
          mem_118 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h77 == io_addr) begin // @[Ram.scala 19:35]
          mem_119 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h78 == io_addr) begin // @[Ram.scala 19:35]
          mem_120 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h79 == io_addr) begin // @[Ram.scala 19:35]
          mem_121 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h7a == io_addr) begin // @[Ram.scala 19:35]
          mem_122 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h7b == io_addr) begin // @[Ram.scala 19:35]
          mem_123 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h7c == io_addr) begin // @[Ram.scala 19:35]
          mem_124 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h7d == io_addr) begin // @[Ram.scala 19:35]
          mem_125 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h7e == io_addr) begin // @[Ram.scala 19:35]
          mem_126 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (7'h7f == io_addr) begin // @[Ram.scala 19:35]
          mem_127 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  mem_0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  mem_1 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  mem_2 = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  mem_3 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  mem_4 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  mem_5 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  mem_6 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  mem_7 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  mem_8 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  mem_9 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  mem_10 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  mem_11 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  mem_12 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  mem_13 = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  mem_14 = _RAND_14[127:0];
  _RAND_15 = {4{`RANDOM}};
  mem_15 = _RAND_15[127:0];
  _RAND_16 = {4{`RANDOM}};
  mem_16 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  mem_17 = _RAND_17[127:0];
  _RAND_18 = {4{`RANDOM}};
  mem_18 = _RAND_18[127:0];
  _RAND_19 = {4{`RANDOM}};
  mem_19 = _RAND_19[127:0];
  _RAND_20 = {4{`RANDOM}};
  mem_20 = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  mem_21 = _RAND_21[127:0];
  _RAND_22 = {4{`RANDOM}};
  mem_22 = _RAND_22[127:0];
  _RAND_23 = {4{`RANDOM}};
  mem_23 = _RAND_23[127:0];
  _RAND_24 = {4{`RANDOM}};
  mem_24 = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  mem_25 = _RAND_25[127:0];
  _RAND_26 = {4{`RANDOM}};
  mem_26 = _RAND_26[127:0];
  _RAND_27 = {4{`RANDOM}};
  mem_27 = _RAND_27[127:0];
  _RAND_28 = {4{`RANDOM}};
  mem_28 = _RAND_28[127:0];
  _RAND_29 = {4{`RANDOM}};
  mem_29 = _RAND_29[127:0];
  _RAND_30 = {4{`RANDOM}};
  mem_30 = _RAND_30[127:0];
  _RAND_31 = {4{`RANDOM}};
  mem_31 = _RAND_31[127:0];
  _RAND_32 = {4{`RANDOM}};
  mem_32 = _RAND_32[127:0];
  _RAND_33 = {4{`RANDOM}};
  mem_33 = _RAND_33[127:0];
  _RAND_34 = {4{`RANDOM}};
  mem_34 = _RAND_34[127:0];
  _RAND_35 = {4{`RANDOM}};
  mem_35 = _RAND_35[127:0];
  _RAND_36 = {4{`RANDOM}};
  mem_36 = _RAND_36[127:0];
  _RAND_37 = {4{`RANDOM}};
  mem_37 = _RAND_37[127:0];
  _RAND_38 = {4{`RANDOM}};
  mem_38 = _RAND_38[127:0];
  _RAND_39 = {4{`RANDOM}};
  mem_39 = _RAND_39[127:0];
  _RAND_40 = {4{`RANDOM}};
  mem_40 = _RAND_40[127:0];
  _RAND_41 = {4{`RANDOM}};
  mem_41 = _RAND_41[127:0];
  _RAND_42 = {4{`RANDOM}};
  mem_42 = _RAND_42[127:0];
  _RAND_43 = {4{`RANDOM}};
  mem_43 = _RAND_43[127:0];
  _RAND_44 = {4{`RANDOM}};
  mem_44 = _RAND_44[127:0];
  _RAND_45 = {4{`RANDOM}};
  mem_45 = _RAND_45[127:0];
  _RAND_46 = {4{`RANDOM}};
  mem_46 = _RAND_46[127:0];
  _RAND_47 = {4{`RANDOM}};
  mem_47 = _RAND_47[127:0];
  _RAND_48 = {4{`RANDOM}};
  mem_48 = _RAND_48[127:0];
  _RAND_49 = {4{`RANDOM}};
  mem_49 = _RAND_49[127:0];
  _RAND_50 = {4{`RANDOM}};
  mem_50 = _RAND_50[127:0];
  _RAND_51 = {4{`RANDOM}};
  mem_51 = _RAND_51[127:0];
  _RAND_52 = {4{`RANDOM}};
  mem_52 = _RAND_52[127:0];
  _RAND_53 = {4{`RANDOM}};
  mem_53 = _RAND_53[127:0];
  _RAND_54 = {4{`RANDOM}};
  mem_54 = _RAND_54[127:0];
  _RAND_55 = {4{`RANDOM}};
  mem_55 = _RAND_55[127:0];
  _RAND_56 = {4{`RANDOM}};
  mem_56 = _RAND_56[127:0];
  _RAND_57 = {4{`RANDOM}};
  mem_57 = _RAND_57[127:0];
  _RAND_58 = {4{`RANDOM}};
  mem_58 = _RAND_58[127:0];
  _RAND_59 = {4{`RANDOM}};
  mem_59 = _RAND_59[127:0];
  _RAND_60 = {4{`RANDOM}};
  mem_60 = _RAND_60[127:0];
  _RAND_61 = {4{`RANDOM}};
  mem_61 = _RAND_61[127:0];
  _RAND_62 = {4{`RANDOM}};
  mem_62 = _RAND_62[127:0];
  _RAND_63 = {4{`RANDOM}};
  mem_63 = _RAND_63[127:0];
  _RAND_64 = {4{`RANDOM}};
  mem_64 = _RAND_64[127:0];
  _RAND_65 = {4{`RANDOM}};
  mem_65 = _RAND_65[127:0];
  _RAND_66 = {4{`RANDOM}};
  mem_66 = _RAND_66[127:0];
  _RAND_67 = {4{`RANDOM}};
  mem_67 = _RAND_67[127:0];
  _RAND_68 = {4{`RANDOM}};
  mem_68 = _RAND_68[127:0];
  _RAND_69 = {4{`RANDOM}};
  mem_69 = _RAND_69[127:0];
  _RAND_70 = {4{`RANDOM}};
  mem_70 = _RAND_70[127:0];
  _RAND_71 = {4{`RANDOM}};
  mem_71 = _RAND_71[127:0];
  _RAND_72 = {4{`RANDOM}};
  mem_72 = _RAND_72[127:0];
  _RAND_73 = {4{`RANDOM}};
  mem_73 = _RAND_73[127:0];
  _RAND_74 = {4{`RANDOM}};
  mem_74 = _RAND_74[127:0];
  _RAND_75 = {4{`RANDOM}};
  mem_75 = _RAND_75[127:0];
  _RAND_76 = {4{`RANDOM}};
  mem_76 = _RAND_76[127:0];
  _RAND_77 = {4{`RANDOM}};
  mem_77 = _RAND_77[127:0];
  _RAND_78 = {4{`RANDOM}};
  mem_78 = _RAND_78[127:0];
  _RAND_79 = {4{`RANDOM}};
  mem_79 = _RAND_79[127:0];
  _RAND_80 = {4{`RANDOM}};
  mem_80 = _RAND_80[127:0];
  _RAND_81 = {4{`RANDOM}};
  mem_81 = _RAND_81[127:0];
  _RAND_82 = {4{`RANDOM}};
  mem_82 = _RAND_82[127:0];
  _RAND_83 = {4{`RANDOM}};
  mem_83 = _RAND_83[127:0];
  _RAND_84 = {4{`RANDOM}};
  mem_84 = _RAND_84[127:0];
  _RAND_85 = {4{`RANDOM}};
  mem_85 = _RAND_85[127:0];
  _RAND_86 = {4{`RANDOM}};
  mem_86 = _RAND_86[127:0];
  _RAND_87 = {4{`RANDOM}};
  mem_87 = _RAND_87[127:0];
  _RAND_88 = {4{`RANDOM}};
  mem_88 = _RAND_88[127:0];
  _RAND_89 = {4{`RANDOM}};
  mem_89 = _RAND_89[127:0];
  _RAND_90 = {4{`RANDOM}};
  mem_90 = _RAND_90[127:0];
  _RAND_91 = {4{`RANDOM}};
  mem_91 = _RAND_91[127:0];
  _RAND_92 = {4{`RANDOM}};
  mem_92 = _RAND_92[127:0];
  _RAND_93 = {4{`RANDOM}};
  mem_93 = _RAND_93[127:0];
  _RAND_94 = {4{`RANDOM}};
  mem_94 = _RAND_94[127:0];
  _RAND_95 = {4{`RANDOM}};
  mem_95 = _RAND_95[127:0];
  _RAND_96 = {4{`RANDOM}};
  mem_96 = _RAND_96[127:0];
  _RAND_97 = {4{`RANDOM}};
  mem_97 = _RAND_97[127:0];
  _RAND_98 = {4{`RANDOM}};
  mem_98 = _RAND_98[127:0];
  _RAND_99 = {4{`RANDOM}};
  mem_99 = _RAND_99[127:0];
  _RAND_100 = {4{`RANDOM}};
  mem_100 = _RAND_100[127:0];
  _RAND_101 = {4{`RANDOM}};
  mem_101 = _RAND_101[127:0];
  _RAND_102 = {4{`RANDOM}};
  mem_102 = _RAND_102[127:0];
  _RAND_103 = {4{`RANDOM}};
  mem_103 = _RAND_103[127:0];
  _RAND_104 = {4{`RANDOM}};
  mem_104 = _RAND_104[127:0];
  _RAND_105 = {4{`RANDOM}};
  mem_105 = _RAND_105[127:0];
  _RAND_106 = {4{`RANDOM}};
  mem_106 = _RAND_106[127:0];
  _RAND_107 = {4{`RANDOM}};
  mem_107 = _RAND_107[127:0];
  _RAND_108 = {4{`RANDOM}};
  mem_108 = _RAND_108[127:0];
  _RAND_109 = {4{`RANDOM}};
  mem_109 = _RAND_109[127:0];
  _RAND_110 = {4{`RANDOM}};
  mem_110 = _RAND_110[127:0];
  _RAND_111 = {4{`RANDOM}};
  mem_111 = _RAND_111[127:0];
  _RAND_112 = {4{`RANDOM}};
  mem_112 = _RAND_112[127:0];
  _RAND_113 = {4{`RANDOM}};
  mem_113 = _RAND_113[127:0];
  _RAND_114 = {4{`RANDOM}};
  mem_114 = _RAND_114[127:0];
  _RAND_115 = {4{`RANDOM}};
  mem_115 = _RAND_115[127:0];
  _RAND_116 = {4{`RANDOM}};
  mem_116 = _RAND_116[127:0];
  _RAND_117 = {4{`RANDOM}};
  mem_117 = _RAND_117[127:0];
  _RAND_118 = {4{`RANDOM}};
  mem_118 = _RAND_118[127:0];
  _RAND_119 = {4{`RANDOM}};
  mem_119 = _RAND_119[127:0];
  _RAND_120 = {4{`RANDOM}};
  mem_120 = _RAND_120[127:0];
  _RAND_121 = {4{`RANDOM}};
  mem_121 = _RAND_121[127:0];
  _RAND_122 = {4{`RANDOM}};
  mem_122 = _RAND_122[127:0];
  _RAND_123 = {4{`RANDOM}};
  mem_123 = _RAND_123[127:0];
  _RAND_124 = {4{`RANDOM}};
  mem_124 = _RAND_124[127:0];
  _RAND_125 = {4{`RANDOM}};
  mem_125 = _RAND_125[127:0];
  _RAND_126 = {4{`RANDOM}};
  mem_126 = _RAND_126[127:0];
  _RAND_127 = {4{`RANDOM}};
  mem_127 = _RAND_127[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
