module RWSmem(
  input          clock,
  input          reset,
  input          io_enable,
  input          io_write,
  input  [9:0]   io_addr,
  input  [255:0] io_dataIn,
  output [255:0] io_dataOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [255:0] _RAND_0;
  reg [255:0] _RAND_1;
  reg [255:0] _RAND_2;
  reg [255:0] _RAND_3;
  reg [255:0] _RAND_4;
  reg [255:0] _RAND_5;
  reg [255:0] _RAND_6;
  reg [255:0] _RAND_7;
  reg [255:0] _RAND_8;
  reg [255:0] _RAND_9;
  reg [255:0] _RAND_10;
  reg [255:0] _RAND_11;
  reg [255:0] _RAND_12;
  reg [255:0] _RAND_13;
  reg [255:0] _RAND_14;
  reg [255:0] _RAND_15;
  reg [255:0] _RAND_16;
  reg [255:0] _RAND_17;
  reg [255:0] _RAND_18;
  reg [255:0] _RAND_19;
  reg [255:0] _RAND_20;
  reg [255:0] _RAND_21;
  reg [255:0] _RAND_22;
  reg [255:0] _RAND_23;
  reg [255:0] _RAND_24;
  reg [255:0] _RAND_25;
  reg [255:0] _RAND_26;
  reg [255:0] _RAND_27;
  reg [255:0] _RAND_28;
  reg [255:0] _RAND_29;
  reg [255:0] _RAND_30;
  reg [255:0] _RAND_31;
  reg [255:0] _RAND_32;
  reg [255:0] _RAND_33;
  reg [255:0] _RAND_34;
  reg [255:0] _RAND_35;
  reg [255:0] _RAND_36;
  reg [255:0] _RAND_37;
  reg [255:0] _RAND_38;
  reg [255:0] _RAND_39;
  reg [255:0] _RAND_40;
  reg [255:0] _RAND_41;
  reg [255:0] _RAND_42;
  reg [255:0] _RAND_43;
  reg [255:0] _RAND_44;
  reg [255:0] _RAND_45;
  reg [255:0] _RAND_46;
  reg [255:0] _RAND_47;
  reg [255:0] _RAND_48;
  reg [255:0] _RAND_49;
  reg [255:0] _RAND_50;
  reg [255:0] _RAND_51;
  reg [255:0] _RAND_52;
  reg [255:0] _RAND_53;
  reg [255:0] _RAND_54;
  reg [255:0] _RAND_55;
  reg [255:0] _RAND_56;
  reg [255:0] _RAND_57;
  reg [255:0] _RAND_58;
  reg [255:0] _RAND_59;
  reg [255:0] _RAND_60;
  reg [255:0] _RAND_61;
  reg [255:0] _RAND_62;
  reg [255:0] _RAND_63;
  reg [255:0] _RAND_64;
  reg [255:0] _RAND_65;
  reg [255:0] _RAND_66;
  reg [255:0] _RAND_67;
  reg [255:0] _RAND_68;
  reg [255:0] _RAND_69;
  reg [255:0] _RAND_70;
  reg [255:0] _RAND_71;
  reg [255:0] _RAND_72;
  reg [255:0] _RAND_73;
  reg [255:0] _RAND_74;
  reg [255:0] _RAND_75;
  reg [255:0] _RAND_76;
  reg [255:0] _RAND_77;
  reg [255:0] _RAND_78;
  reg [255:0] _RAND_79;
  reg [255:0] _RAND_80;
  reg [255:0] _RAND_81;
  reg [255:0] _RAND_82;
  reg [255:0] _RAND_83;
  reg [255:0] _RAND_84;
  reg [255:0] _RAND_85;
  reg [255:0] _RAND_86;
  reg [255:0] _RAND_87;
  reg [255:0] _RAND_88;
  reg [255:0] _RAND_89;
  reg [255:0] _RAND_90;
  reg [255:0] _RAND_91;
  reg [255:0] _RAND_92;
  reg [255:0] _RAND_93;
  reg [255:0] _RAND_94;
  reg [255:0] _RAND_95;
  reg [255:0] _RAND_96;
  reg [255:0] _RAND_97;
  reg [255:0] _RAND_98;
  reg [255:0] _RAND_99;
  reg [255:0] _RAND_100;
  reg [255:0] _RAND_101;
  reg [255:0] _RAND_102;
  reg [255:0] _RAND_103;
  reg [255:0] _RAND_104;
  reg [255:0] _RAND_105;
  reg [255:0] _RAND_106;
  reg [255:0] _RAND_107;
  reg [255:0] _RAND_108;
  reg [255:0] _RAND_109;
  reg [255:0] _RAND_110;
  reg [255:0] _RAND_111;
  reg [255:0] _RAND_112;
  reg [255:0] _RAND_113;
  reg [255:0] _RAND_114;
  reg [255:0] _RAND_115;
  reg [255:0] _RAND_116;
  reg [255:0] _RAND_117;
  reg [255:0] _RAND_118;
  reg [255:0] _RAND_119;
  reg [255:0] _RAND_120;
  reg [255:0] _RAND_121;
  reg [255:0] _RAND_122;
  reg [255:0] _RAND_123;
  reg [255:0] _RAND_124;
  reg [255:0] _RAND_125;
  reg [255:0] _RAND_126;
  reg [255:0] _RAND_127;
  reg [255:0] _RAND_128;
  reg [255:0] _RAND_129;
  reg [255:0] _RAND_130;
  reg [255:0] _RAND_131;
  reg [255:0] _RAND_132;
  reg [255:0] _RAND_133;
  reg [255:0] _RAND_134;
  reg [255:0] _RAND_135;
  reg [255:0] _RAND_136;
  reg [255:0] _RAND_137;
  reg [255:0] _RAND_138;
  reg [255:0] _RAND_139;
  reg [255:0] _RAND_140;
  reg [255:0] _RAND_141;
  reg [255:0] _RAND_142;
  reg [255:0] _RAND_143;
  reg [255:0] _RAND_144;
  reg [255:0] _RAND_145;
  reg [255:0] _RAND_146;
  reg [255:0] _RAND_147;
  reg [255:0] _RAND_148;
  reg [255:0] _RAND_149;
  reg [255:0] _RAND_150;
  reg [255:0] _RAND_151;
  reg [255:0] _RAND_152;
  reg [255:0] _RAND_153;
  reg [255:0] _RAND_154;
  reg [255:0] _RAND_155;
  reg [255:0] _RAND_156;
  reg [255:0] _RAND_157;
  reg [255:0] _RAND_158;
  reg [255:0] _RAND_159;
  reg [255:0] _RAND_160;
  reg [255:0] _RAND_161;
  reg [255:0] _RAND_162;
  reg [255:0] _RAND_163;
  reg [255:0] _RAND_164;
  reg [255:0] _RAND_165;
  reg [255:0] _RAND_166;
  reg [255:0] _RAND_167;
  reg [255:0] _RAND_168;
  reg [255:0] _RAND_169;
  reg [255:0] _RAND_170;
  reg [255:0] _RAND_171;
  reg [255:0] _RAND_172;
  reg [255:0] _RAND_173;
  reg [255:0] _RAND_174;
  reg [255:0] _RAND_175;
  reg [255:0] _RAND_176;
  reg [255:0] _RAND_177;
  reg [255:0] _RAND_178;
  reg [255:0] _RAND_179;
  reg [255:0] _RAND_180;
  reg [255:0] _RAND_181;
  reg [255:0] _RAND_182;
  reg [255:0] _RAND_183;
  reg [255:0] _RAND_184;
  reg [255:0] _RAND_185;
  reg [255:0] _RAND_186;
  reg [255:0] _RAND_187;
  reg [255:0] _RAND_188;
  reg [255:0] _RAND_189;
  reg [255:0] _RAND_190;
  reg [255:0] _RAND_191;
  reg [255:0] _RAND_192;
  reg [255:0] _RAND_193;
  reg [255:0] _RAND_194;
  reg [255:0] _RAND_195;
  reg [255:0] _RAND_196;
  reg [255:0] _RAND_197;
  reg [255:0] _RAND_198;
  reg [255:0] _RAND_199;
  reg [255:0] _RAND_200;
  reg [255:0] _RAND_201;
  reg [255:0] _RAND_202;
  reg [255:0] _RAND_203;
  reg [255:0] _RAND_204;
  reg [255:0] _RAND_205;
  reg [255:0] _RAND_206;
  reg [255:0] _RAND_207;
  reg [255:0] _RAND_208;
  reg [255:0] _RAND_209;
  reg [255:0] _RAND_210;
  reg [255:0] _RAND_211;
  reg [255:0] _RAND_212;
  reg [255:0] _RAND_213;
  reg [255:0] _RAND_214;
  reg [255:0] _RAND_215;
  reg [255:0] _RAND_216;
  reg [255:0] _RAND_217;
  reg [255:0] _RAND_218;
  reg [255:0] _RAND_219;
  reg [255:0] _RAND_220;
  reg [255:0] _RAND_221;
  reg [255:0] _RAND_222;
  reg [255:0] _RAND_223;
  reg [255:0] _RAND_224;
  reg [255:0] _RAND_225;
  reg [255:0] _RAND_226;
  reg [255:0] _RAND_227;
  reg [255:0] _RAND_228;
  reg [255:0] _RAND_229;
  reg [255:0] _RAND_230;
  reg [255:0] _RAND_231;
  reg [255:0] _RAND_232;
  reg [255:0] _RAND_233;
  reg [255:0] _RAND_234;
  reg [255:0] _RAND_235;
  reg [255:0] _RAND_236;
  reg [255:0] _RAND_237;
  reg [255:0] _RAND_238;
  reg [255:0] _RAND_239;
  reg [255:0] _RAND_240;
  reg [255:0] _RAND_241;
  reg [255:0] _RAND_242;
  reg [255:0] _RAND_243;
  reg [255:0] _RAND_244;
  reg [255:0] _RAND_245;
  reg [255:0] _RAND_246;
  reg [255:0] _RAND_247;
  reg [255:0] _RAND_248;
  reg [255:0] _RAND_249;
  reg [255:0] _RAND_250;
  reg [255:0] _RAND_251;
  reg [255:0] _RAND_252;
  reg [255:0] _RAND_253;
  reg [255:0] _RAND_254;
  reg [255:0] _RAND_255;
  reg [255:0] _RAND_256;
  reg [255:0] _RAND_257;
  reg [255:0] _RAND_258;
  reg [255:0] _RAND_259;
  reg [255:0] _RAND_260;
  reg [255:0] _RAND_261;
  reg [255:0] _RAND_262;
  reg [255:0] _RAND_263;
  reg [255:0] _RAND_264;
  reg [255:0] _RAND_265;
  reg [255:0] _RAND_266;
  reg [255:0] _RAND_267;
  reg [255:0] _RAND_268;
  reg [255:0] _RAND_269;
  reg [255:0] _RAND_270;
  reg [255:0] _RAND_271;
  reg [255:0] _RAND_272;
  reg [255:0] _RAND_273;
  reg [255:0] _RAND_274;
  reg [255:0] _RAND_275;
  reg [255:0] _RAND_276;
  reg [255:0] _RAND_277;
  reg [255:0] _RAND_278;
  reg [255:0] _RAND_279;
  reg [255:0] _RAND_280;
  reg [255:0] _RAND_281;
  reg [255:0] _RAND_282;
  reg [255:0] _RAND_283;
  reg [255:0] _RAND_284;
  reg [255:0] _RAND_285;
  reg [255:0] _RAND_286;
  reg [255:0] _RAND_287;
  reg [255:0] _RAND_288;
  reg [255:0] _RAND_289;
  reg [255:0] _RAND_290;
  reg [255:0] _RAND_291;
  reg [255:0] _RAND_292;
  reg [255:0] _RAND_293;
  reg [255:0] _RAND_294;
  reg [255:0] _RAND_295;
  reg [255:0] _RAND_296;
  reg [255:0] _RAND_297;
  reg [255:0] _RAND_298;
  reg [255:0] _RAND_299;
  reg [255:0] _RAND_300;
  reg [255:0] _RAND_301;
  reg [255:0] _RAND_302;
  reg [255:0] _RAND_303;
  reg [255:0] _RAND_304;
  reg [255:0] _RAND_305;
  reg [255:0] _RAND_306;
  reg [255:0] _RAND_307;
  reg [255:0] _RAND_308;
  reg [255:0] _RAND_309;
  reg [255:0] _RAND_310;
  reg [255:0] _RAND_311;
  reg [255:0] _RAND_312;
  reg [255:0] _RAND_313;
  reg [255:0] _RAND_314;
  reg [255:0] _RAND_315;
  reg [255:0] _RAND_316;
  reg [255:0] _RAND_317;
  reg [255:0] _RAND_318;
  reg [255:0] _RAND_319;
  reg [255:0] _RAND_320;
  reg [255:0] _RAND_321;
  reg [255:0] _RAND_322;
  reg [255:0] _RAND_323;
  reg [255:0] _RAND_324;
  reg [255:0] _RAND_325;
  reg [255:0] _RAND_326;
  reg [255:0] _RAND_327;
  reg [255:0] _RAND_328;
  reg [255:0] _RAND_329;
  reg [255:0] _RAND_330;
  reg [255:0] _RAND_331;
  reg [255:0] _RAND_332;
  reg [255:0] _RAND_333;
  reg [255:0] _RAND_334;
  reg [255:0] _RAND_335;
  reg [255:0] _RAND_336;
  reg [255:0] _RAND_337;
  reg [255:0] _RAND_338;
  reg [255:0] _RAND_339;
  reg [255:0] _RAND_340;
  reg [255:0] _RAND_341;
  reg [255:0] _RAND_342;
  reg [255:0] _RAND_343;
  reg [255:0] _RAND_344;
  reg [255:0] _RAND_345;
  reg [255:0] _RAND_346;
  reg [255:0] _RAND_347;
  reg [255:0] _RAND_348;
  reg [255:0] _RAND_349;
  reg [255:0] _RAND_350;
  reg [255:0] _RAND_351;
  reg [255:0] _RAND_352;
  reg [255:0] _RAND_353;
  reg [255:0] _RAND_354;
  reg [255:0] _RAND_355;
  reg [255:0] _RAND_356;
  reg [255:0] _RAND_357;
  reg [255:0] _RAND_358;
  reg [255:0] _RAND_359;
  reg [255:0] _RAND_360;
  reg [255:0] _RAND_361;
  reg [255:0] _RAND_362;
  reg [255:0] _RAND_363;
  reg [255:0] _RAND_364;
  reg [255:0] _RAND_365;
  reg [255:0] _RAND_366;
  reg [255:0] _RAND_367;
  reg [255:0] _RAND_368;
  reg [255:0] _RAND_369;
  reg [255:0] _RAND_370;
  reg [255:0] _RAND_371;
  reg [255:0] _RAND_372;
  reg [255:0] _RAND_373;
  reg [255:0] _RAND_374;
  reg [255:0] _RAND_375;
  reg [255:0] _RAND_376;
  reg [255:0] _RAND_377;
  reg [255:0] _RAND_378;
  reg [255:0] _RAND_379;
  reg [255:0] _RAND_380;
  reg [255:0] _RAND_381;
  reg [255:0] _RAND_382;
  reg [255:0] _RAND_383;
  reg [255:0] _RAND_384;
  reg [255:0] _RAND_385;
  reg [255:0] _RAND_386;
  reg [255:0] _RAND_387;
  reg [255:0] _RAND_388;
  reg [255:0] _RAND_389;
  reg [255:0] _RAND_390;
  reg [255:0] _RAND_391;
  reg [255:0] _RAND_392;
  reg [255:0] _RAND_393;
  reg [255:0] _RAND_394;
  reg [255:0] _RAND_395;
  reg [255:0] _RAND_396;
  reg [255:0] _RAND_397;
  reg [255:0] _RAND_398;
  reg [255:0] _RAND_399;
  reg [255:0] _RAND_400;
  reg [255:0] _RAND_401;
  reg [255:0] _RAND_402;
  reg [255:0] _RAND_403;
  reg [255:0] _RAND_404;
  reg [255:0] _RAND_405;
  reg [255:0] _RAND_406;
  reg [255:0] _RAND_407;
  reg [255:0] _RAND_408;
  reg [255:0] _RAND_409;
  reg [255:0] _RAND_410;
  reg [255:0] _RAND_411;
  reg [255:0] _RAND_412;
  reg [255:0] _RAND_413;
  reg [255:0] _RAND_414;
  reg [255:0] _RAND_415;
  reg [255:0] _RAND_416;
  reg [255:0] _RAND_417;
  reg [255:0] _RAND_418;
  reg [255:0] _RAND_419;
  reg [255:0] _RAND_420;
  reg [255:0] _RAND_421;
  reg [255:0] _RAND_422;
  reg [255:0] _RAND_423;
  reg [255:0] _RAND_424;
  reg [255:0] _RAND_425;
  reg [255:0] _RAND_426;
  reg [255:0] _RAND_427;
  reg [255:0] _RAND_428;
  reg [255:0] _RAND_429;
  reg [255:0] _RAND_430;
  reg [255:0] _RAND_431;
  reg [255:0] _RAND_432;
  reg [255:0] _RAND_433;
  reg [255:0] _RAND_434;
  reg [255:0] _RAND_435;
  reg [255:0] _RAND_436;
  reg [255:0] _RAND_437;
  reg [255:0] _RAND_438;
  reg [255:0] _RAND_439;
  reg [255:0] _RAND_440;
  reg [255:0] _RAND_441;
  reg [255:0] _RAND_442;
  reg [255:0] _RAND_443;
  reg [255:0] _RAND_444;
  reg [255:0] _RAND_445;
  reg [255:0] _RAND_446;
  reg [255:0] _RAND_447;
  reg [255:0] _RAND_448;
  reg [255:0] _RAND_449;
  reg [255:0] _RAND_450;
  reg [255:0] _RAND_451;
  reg [255:0] _RAND_452;
  reg [255:0] _RAND_453;
  reg [255:0] _RAND_454;
  reg [255:0] _RAND_455;
  reg [255:0] _RAND_456;
  reg [255:0] _RAND_457;
  reg [255:0] _RAND_458;
  reg [255:0] _RAND_459;
  reg [255:0] _RAND_460;
  reg [255:0] _RAND_461;
  reg [255:0] _RAND_462;
  reg [255:0] _RAND_463;
  reg [255:0] _RAND_464;
  reg [255:0] _RAND_465;
  reg [255:0] _RAND_466;
  reg [255:0] _RAND_467;
  reg [255:0] _RAND_468;
  reg [255:0] _RAND_469;
  reg [255:0] _RAND_470;
  reg [255:0] _RAND_471;
  reg [255:0] _RAND_472;
  reg [255:0] _RAND_473;
  reg [255:0] _RAND_474;
  reg [255:0] _RAND_475;
  reg [255:0] _RAND_476;
  reg [255:0] _RAND_477;
  reg [255:0] _RAND_478;
  reg [255:0] _RAND_479;
  reg [255:0] _RAND_480;
  reg [255:0] _RAND_481;
  reg [255:0] _RAND_482;
  reg [255:0] _RAND_483;
  reg [255:0] _RAND_484;
  reg [255:0] _RAND_485;
  reg [255:0] _RAND_486;
  reg [255:0] _RAND_487;
  reg [255:0] _RAND_488;
  reg [255:0] _RAND_489;
  reg [255:0] _RAND_490;
  reg [255:0] _RAND_491;
  reg [255:0] _RAND_492;
  reg [255:0] _RAND_493;
  reg [255:0] _RAND_494;
  reg [255:0] _RAND_495;
  reg [255:0] _RAND_496;
  reg [255:0] _RAND_497;
  reg [255:0] _RAND_498;
  reg [255:0] _RAND_499;
  reg [255:0] _RAND_500;
  reg [255:0] _RAND_501;
  reg [255:0] _RAND_502;
  reg [255:0] _RAND_503;
  reg [255:0] _RAND_504;
  reg [255:0] _RAND_505;
  reg [255:0] _RAND_506;
  reg [255:0] _RAND_507;
  reg [255:0] _RAND_508;
  reg [255:0] _RAND_509;
  reg [255:0] _RAND_510;
  reg [255:0] _RAND_511;
  reg [255:0] _RAND_512;
  reg [255:0] _RAND_513;
  reg [255:0] _RAND_514;
  reg [255:0] _RAND_515;
  reg [255:0] _RAND_516;
  reg [255:0] _RAND_517;
  reg [255:0] _RAND_518;
  reg [255:0] _RAND_519;
  reg [255:0] _RAND_520;
  reg [255:0] _RAND_521;
  reg [255:0] _RAND_522;
  reg [255:0] _RAND_523;
  reg [255:0] _RAND_524;
  reg [255:0] _RAND_525;
  reg [255:0] _RAND_526;
  reg [255:0] _RAND_527;
  reg [255:0] _RAND_528;
  reg [255:0] _RAND_529;
  reg [255:0] _RAND_530;
  reg [255:0] _RAND_531;
  reg [255:0] _RAND_532;
  reg [255:0] _RAND_533;
  reg [255:0] _RAND_534;
  reg [255:0] _RAND_535;
  reg [255:0] _RAND_536;
  reg [255:0] _RAND_537;
  reg [255:0] _RAND_538;
  reg [255:0] _RAND_539;
  reg [255:0] _RAND_540;
  reg [255:0] _RAND_541;
  reg [255:0] _RAND_542;
  reg [255:0] _RAND_543;
  reg [255:0] _RAND_544;
  reg [255:0] _RAND_545;
  reg [255:0] _RAND_546;
  reg [255:0] _RAND_547;
  reg [255:0] _RAND_548;
  reg [255:0] _RAND_549;
  reg [255:0] _RAND_550;
  reg [255:0] _RAND_551;
  reg [255:0] _RAND_552;
  reg [255:0] _RAND_553;
  reg [255:0] _RAND_554;
  reg [255:0] _RAND_555;
  reg [255:0] _RAND_556;
  reg [255:0] _RAND_557;
  reg [255:0] _RAND_558;
  reg [255:0] _RAND_559;
  reg [255:0] _RAND_560;
  reg [255:0] _RAND_561;
  reg [255:0] _RAND_562;
  reg [255:0] _RAND_563;
  reg [255:0] _RAND_564;
  reg [255:0] _RAND_565;
  reg [255:0] _RAND_566;
  reg [255:0] _RAND_567;
  reg [255:0] _RAND_568;
  reg [255:0] _RAND_569;
  reg [255:0] _RAND_570;
  reg [255:0] _RAND_571;
  reg [255:0] _RAND_572;
  reg [255:0] _RAND_573;
  reg [255:0] _RAND_574;
  reg [255:0] _RAND_575;
  reg [255:0] _RAND_576;
  reg [255:0] _RAND_577;
  reg [255:0] _RAND_578;
  reg [255:0] _RAND_579;
  reg [255:0] _RAND_580;
  reg [255:0] _RAND_581;
  reg [255:0] _RAND_582;
  reg [255:0] _RAND_583;
  reg [255:0] _RAND_584;
  reg [255:0] _RAND_585;
  reg [255:0] _RAND_586;
  reg [255:0] _RAND_587;
  reg [255:0] _RAND_588;
  reg [255:0] _RAND_589;
  reg [255:0] _RAND_590;
  reg [255:0] _RAND_591;
  reg [255:0] _RAND_592;
  reg [255:0] _RAND_593;
  reg [255:0] _RAND_594;
  reg [255:0] _RAND_595;
  reg [255:0] _RAND_596;
  reg [255:0] _RAND_597;
  reg [255:0] _RAND_598;
  reg [255:0] _RAND_599;
  reg [255:0] _RAND_600;
  reg [255:0] _RAND_601;
  reg [255:0] _RAND_602;
  reg [255:0] _RAND_603;
  reg [255:0] _RAND_604;
  reg [255:0] _RAND_605;
  reg [255:0] _RAND_606;
  reg [255:0] _RAND_607;
  reg [255:0] _RAND_608;
  reg [255:0] _RAND_609;
  reg [255:0] _RAND_610;
  reg [255:0] _RAND_611;
  reg [255:0] _RAND_612;
  reg [255:0] _RAND_613;
  reg [255:0] _RAND_614;
  reg [255:0] _RAND_615;
  reg [255:0] _RAND_616;
  reg [255:0] _RAND_617;
  reg [255:0] _RAND_618;
  reg [255:0] _RAND_619;
  reg [255:0] _RAND_620;
  reg [255:0] _RAND_621;
  reg [255:0] _RAND_622;
  reg [255:0] _RAND_623;
  reg [255:0] _RAND_624;
  reg [255:0] _RAND_625;
  reg [255:0] _RAND_626;
  reg [255:0] _RAND_627;
  reg [255:0] _RAND_628;
  reg [255:0] _RAND_629;
  reg [255:0] _RAND_630;
  reg [255:0] _RAND_631;
  reg [255:0] _RAND_632;
  reg [255:0] _RAND_633;
  reg [255:0] _RAND_634;
  reg [255:0] _RAND_635;
  reg [255:0] _RAND_636;
  reg [255:0] _RAND_637;
  reg [255:0] _RAND_638;
  reg [255:0] _RAND_639;
  reg [255:0] _RAND_640;
  reg [255:0] _RAND_641;
  reg [255:0] _RAND_642;
  reg [255:0] _RAND_643;
  reg [255:0] _RAND_644;
  reg [255:0] _RAND_645;
  reg [255:0] _RAND_646;
  reg [255:0] _RAND_647;
  reg [255:0] _RAND_648;
  reg [255:0] _RAND_649;
  reg [255:0] _RAND_650;
  reg [255:0] _RAND_651;
  reg [255:0] _RAND_652;
  reg [255:0] _RAND_653;
  reg [255:0] _RAND_654;
  reg [255:0] _RAND_655;
  reg [255:0] _RAND_656;
  reg [255:0] _RAND_657;
  reg [255:0] _RAND_658;
  reg [255:0] _RAND_659;
  reg [255:0] _RAND_660;
  reg [255:0] _RAND_661;
  reg [255:0] _RAND_662;
  reg [255:0] _RAND_663;
  reg [255:0] _RAND_664;
  reg [255:0] _RAND_665;
  reg [255:0] _RAND_666;
  reg [255:0] _RAND_667;
  reg [255:0] _RAND_668;
  reg [255:0] _RAND_669;
  reg [255:0] _RAND_670;
  reg [255:0] _RAND_671;
  reg [255:0] _RAND_672;
  reg [255:0] _RAND_673;
  reg [255:0] _RAND_674;
  reg [255:0] _RAND_675;
  reg [255:0] _RAND_676;
  reg [255:0] _RAND_677;
  reg [255:0] _RAND_678;
  reg [255:0] _RAND_679;
  reg [255:0] _RAND_680;
  reg [255:0] _RAND_681;
  reg [255:0] _RAND_682;
  reg [255:0] _RAND_683;
  reg [255:0] _RAND_684;
  reg [255:0] _RAND_685;
  reg [255:0] _RAND_686;
  reg [255:0] _RAND_687;
  reg [255:0] _RAND_688;
  reg [255:0] _RAND_689;
  reg [255:0] _RAND_690;
  reg [255:0] _RAND_691;
  reg [255:0] _RAND_692;
  reg [255:0] _RAND_693;
  reg [255:0] _RAND_694;
  reg [255:0] _RAND_695;
  reg [255:0] _RAND_696;
  reg [255:0] _RAND_697;
  reg [255:0] _RAND_698;
  reg [255:0] _RAND_699;
  reg [255:0] _RAND_700;
  reg [255:0] _RAND_701;
  reg [255:0] _RAND_702;
  reg [255:0] _RAND_703;
  reg [255:0] _RAND_704;
  reg [255:0] _RAND_705;
  reg [255:0] _RAND_706;
  reg [255:0] _RAND_707;
  reg [255:0] _RAND_708;
  reg [255:0] _RAND_709;
  reg [255:0] _RAND_710;
  reg [255:0] _RAND_711;
  reg [255:0] _RAND_712;
  reg [255:0] _RAND_713;
  reg [255:0] _RAND_714;
  reg [255:0] _RAND_715;
  reg [255:0] _RAND_716;
  reg [255:0] _RAND_717;
  reg [255:0] _RAND_718;
  reg [255:0] _RAND_719;
  reg [255:0] _RAND_720;
  reg [255:0] _RAND_721;
  reg [255:0] _RAND_722;
  reg [255:0] _RAND_723;
  reg [255:0] _RAND_724;
  reg [255:0] _RAND_725;
  reg [255:0] _RAND_726;
  reg [255:0] _RAND_727;
  reg [255:0] _RAND_728;
  reg [255:0] _RAND_729;
  reg [255:0] _RAND_730;
  reg [255:0] _RAND_731;
  reg [255:0] _RAND_732;
  reg [255:0] _RAND_733;
  reg [255:0] _RAND_734;
  reg [255:0] _RAND_735;
  reg [255:0] _RAND_736;
  reg [255:0] _RAND_737;
  reg [255:0] _RAND_738;
  reg [255:0] _RAND_739;
  reg [255:0] _RAND_740;
  reg [255:0] _RAND_741;
  reg [255:0] _RAND_742;
  reg [255:0] _RAND_743;
  reg [255:0] _RAND_744;
  reg [255:0] _RAND_745;
  reg [255:0] _RAND_746;
  reg [255:0] _RAND_747;
  reg [255:0] _RAND_748;
  reg [255:0] _RAND_749;
  reg [255:0] _RAND_750;
  reg [255:0] _RAND_751;
  reg [255:0] _RAND_752;
  reg [255:0] _RAND_753;
  reg [255:0] _RAND_754;
  reg [255:0] _RAND_755;
  reg [255:0] _RAND_756;
  reg [255:0] _RAND_757;
  reg [255:0] _RAND_758;
  reg [255:0] _RAND_759;
  reg [255:0] _RAND_760;
  reg [255:0] _RAND_761;
  reg [255:0] _RAND_762;
  reg [255:0] _RAND_763;
  reg [255:0] _RAND_764;
  reg [255:0] _RAND_765;
  reg [255:0] _RAND_766;
  reg [255:0] _RAND_767;
  reg [255:0] _RAND_768;
  reg [255:0] _RAND_769;
  reg [255:0] _RAND_770;
  reg [255:0] _RAND_771;
  reg [255:0] _RAND_772;
  reg [255:0] _RAND_773;
  reg [255:0] _RAND_774;
  reg [255:0] _RAND_775;
  reg [255:0] _RAND_776;
  reg [255:0] _RAND_777;
  reg [255:0] _RAND_778;
  reg [255:0] _RAND_779;
  reg [255:0] _RAND_780;
  reg [255:0] _RAND_781;
  reg [255:0] _RAND_782;
  reg [255:0] _RAND_783;
  reg [255:0] _RAND_784;
  reg [255:0] _RAND_785;
  reg [255:0] _RAND_786;
  reg [255:0] _RAND_787;
  reg [255:0] _RAND_788;
  reg [255:0] _RAND_789;
  reg [255:0] _RAND_790;
  reg [255:0] _RAND_791;
  reg [255:0] _RAND_792;
  reg [255:0] _RAND_793;
  reg [255:0] _RAND_794;
  reg [255:0] _RAND_795;
  reg [255:0] _RAND_796;
  reg [255:0] _RAND_797;
  reg [255:0] _RAND_798;
  reg [255:0] _RAND_799;
  reg [255:0] _RAND_800;
  reg [255:0] _RAND_801;
  reg [255:0] _RAND_802;
  reg [255:0] _RAND_803;
  reg [255:0] _RAND_804;
  reg [255:0] _RAND_805;
  reg [255:0] _RAND_806;
  reg [255:0] _RAND_807;
  reg [255:0] _RAND_808;
  reg [255:0] _RAND_809;
  reg [255:0] _RAND_810;
  reg [255:0] _RAND_811;
  reg [255:0] _RAND_812;
  reg [255:0] _RAND_813;
  reg [255:0] _RAND_814;
  reg [255:0] _RAND_815;
  reg [255:0] _RAND_816;
  reg [255:0] _RAND_817;
  reg [255:0] _RAND_818;
  reg [255:0] _RAND_819;
  reg [255:0] _RAND_820;
  reg [255:0] _RAND_821;
  reg [255:0] _RAND_822;
  reg [255:0] _RAND_823;
  reg [255:0] _RAND_824;
  reg [255:0] _RAND_825;
  reg [255:0] _RAND_826;
  reg [255:0] _RAND_827;
  reg [255:0] _RAND_828;
  reg [255:0] _RAND_829;
  reg [255:0] _RAND_830;
  reg [255:0] _RAND_831;
  reg [255:0] _RAND_832;
  reg [255:0] _RAND_833;
  reg [255:0] _RAND_834;
  reg [255:0] _RAND_835;
  reg [255:0] _RAND_836;
  reg [255:0] _RAND_837;
  reg [255:0] _RAND_838;
  reg [255:0] _RAND_839;
  reg [255:0] _RAND_840;
  reg [255:0] _RAND_841;
  reg [255:0] _RAND_842;
  reg [255:0] _RAND_843;
  reg [255:0] _RAND_844;
  reg [255:0] _RAND_845;
  reg [255:0] _RAND_846;
  reg [255:0] _RAND_847;
  reg [255:0] _RAND_848;
  reg [255:0] _RAND_849;
  reg [255:0] _RAND_850;
  reg [255:0] _RAND_851;
  reg [255:0] _RAND_852;
  reg [255:0] _RAND_853;
  reg [255:0] _RAND_854;
  reg [255:0] _RAND_855;
  reg [255:0] _RAND_856;
  reg [255:0] _RAND_857;
  reg [255:0] _RAND_858;
  reg [255:0] _RAND_859;
  reg [255:0] _RAND_860;
  reg [255:0] _RAND_861;
  reg [255:0] _RAND_862;
  reg [255:0] _RAND_863;
  reg [255:0] _RAND_864;
  reg [255:0] _RAND_865;
  reg [255:0] _RAND_866;
  reg [255:0] _RAND_867;
  reg [255:0] _RAND_868;
  reg [255:0] _RAND_869;
  reg [255:0] _RAND_870;
  reg [255:0] _RAND_871;
  reg [255:0] _RAND_872;
  reg [255:0] _RAND_873;
  reg [255:0] _RAND_874;
  reg [255:0] _RAND_875;
  reg [255:0] _RAND_876;
  reg [255:0] _RAND_877;
  reg [255:0] _RAND_878;
  reg [255:0] _RAND_879;
  reg [255:0] _RAND_880;
  reg [255:0] _RAND_881;
  reg [255:0] _RAND_882;
  reg [255:0] _RAND_883;
  reg [255:0] _RAND_884;
  reg [255:0] _RAND_885;
  reg [255:0] _RAND_886;
  reg [255:0] _RAND_887;
  reg [255:0] _RAND_888;
  reg [255:0] _RAND_889;
  reg [255:0] _RAND_890;
  reg [255:0] _RAND_891;
  reg [255:0] _RAND_892;
  reg [255:0] _RAND_893;
  reg [255:0] _RAND_894;
  reg [255:0] _RAND_895;
  reg [255:0] _RAND_896;
  reg [255:0] _RAND_897;
  reg [255:0] _RAND_898;
  reg [255:0] _RAND_899;
  reg [255:0] _RAND_900;
  reg [255:0] _RAND_901;
  reg [255:0] _RAND_902;
  reg [255:0] _RAND_903;
  reg [255:0] _RAND_904;
  reg [255:0] _RAND_905;
  reg [255:0] _RAND_906;
  reg [255:0] _RAND_907;
  reg [255:0] _RAND_908;
  reg [255:0] _RAND_909;
  reg [255:0] _RAND_910;
  reg [255:0] _RAND_911;
  reg [255:0] _RAND_912;
  reg [255:0] _RAND_913;
  reg [255:0] _RAND_914;
  reg [255:0] _RAND_915;
  reg [255:0] _RAND_916;
  reg [255:0] _RAND_917;
  reg [255:0] _RAND_918;
  reg [255:0] _RAND_919;
  reg [255:0] _RAND_920;
  reg [255:0] _RAND_921;
  reg [255:0] _RAND_922;
  reg [255:0] _RAND_923;
  reg [255:0] _RAND_924;
  reg [255:0] _RAND_925;
  reg [255:0] _RAND_926;
  reg [255:0] _RAND_927;
  reg [255:0] _RAND_928;
  reg [255:0] _RAND_929;
  reg [255:0] _RAND_930;
  reg [255:0] _RAND_931;
  reg [255:0] _RAND_932;
  reg [255:0] _RAND_933;
  reg [255:0] _RAND_934;
  reg [255:0] _RAND_935;
  reg [255:0] _RAND_936;
  reg [255:0] _RAND_937;
  reg [255:0] _RAND_938;
  reg [255:0] _RAND_939;
  reg [255:0] _RAND_940;
  reg [255:0] _RAND_941;
  reg [255:0] _RAND_942;
  reg [255:0] _RAND_943;
  reg [255:0] _RAND_944;
  reg [255:0] _RAND_945;
  reg [255:0] _RAND_946;
  reg [255:0] _RAND_947;
  reg [255:0] _RAND_948;
  reg [255:0] _RAND_949;
  reg [255:0] _RAND_950;
  reg [255:0] _RAND_951;
  reg [255:0] _RAND_952;
  reg [255:0] _RAND_953;
  reg [255:0] _RAND_954;
  reg [255:0] _RAND_955;
  reg [255:0] _RAND_956;
  reg [255:0] _RAND_957;
  reg [255:0] _RAND_958;
  reg [255:0] _RAND_959;
  reg [255:0] _RAND_960;
  reg [255:0] _RAND_961;
  reg [255:0] _RAND_962;
  reg [255:0] _RAND_963;
  reg [255:0] _RAND_964;
  reg [255:0] _RAND_965;
  reg [255:0] _RAND_966;
  reg [255:0] _RAND_967;
  reg [255:0] _RAND_968;
  reg [255:0] _RAND_969;
  reg [255:0] _RAND_970;
  reg [255:0] _RAND_971;
  reg [255:0] _RAND_972;
  reg [255:0] _RAND_973;
  reg [255:0] _RAND_974;
  reg [255:0] _RAND_975;
  reg [255:0] _RAND_976;
  reg [255:0] _RAND_977;
  reg [255:0] _RAND_978;
  reg [255:0] _RAND_979;
  reg [255:0] _RAND_980;
  reg [255:0] _RAND_981;
  reg [255:0] _RAND_982;
  reg [255:0] _RAND_983;
  reg [255:0] _RAND_984;
  reg [255:0] _RAND_985;
  reg [255:0] _RAND_986;
  reg [255:0] _RAND_987;
  reg [255:0] _RAND_988;
  reg [255:0] _RAND_989;
  reg [255:0] _RAND_990;
  reg [255:0] _RAND_991;
  reg [255:0] _RAND_992;
  reg [255:0] _RAND_993;
  reg [255:0] _RAND_994;
  reg [255:0] _RAND_995;
  reg [255:0] _RAND_996;
  reg [255:0] _RAND_997;
  reg [255:0] _RAND_998;
  reg [255:0] _RAND_999;
  reg [255:0] _RAND_1000;
  reg [255:0] _RAND_1001;
  reg [255:0] _RAND_1002;
  reg [255:0] _RAND_1003;
  reg [255:0] _RAND_1004;
  reg [255:0] _RAND_1005;
  reg [255:0] _RAND_1006;
  reg [255:0] _RAND_1007;
  reg [255:0] _RAND_1008;
  reg [255:0] _RAND_1009;
  reg [255:0] _RAND_1010;
  reg [255:0] _RAND_1011;
  reg [255:0] _RAND_1012;
  reg [255:0] _RAND_1013;
  reg [255:0] _RAND_1014;
  reg [255:0] _RAND_1015;
  reg [255:0] _RAND_1016;
  reg [255:0] _RAND_1017;
  reg [255:0] _RAND_1018;
  reg [255:0] _RAND_1019;
  reg [255:0] _RAND_1020;
  reg [255:0] _RAND_1021;
  reg [255:0] _RAND_1022;
  reg [255:0] _RAND_1023;
`endif // RANDOMIZE_REG_INIT
  reg [255:0] mem_0; // @[Ram.scala 16:16]
  reg [255:0] mem_1; // @[Ram.scala 16:16]
  reg [255:0] mem_2; // @[Ram.scala 16:16]
  reg [255:0] mem_3; // @[Ram.scala 16:16]
  reg [255:0] mem_4; // @[Ram.scala 16:16]
  reg [255:0] mem_5; // @[Ram.scala 16:16]
  reg [255:0] mem_6; // @[Ram.scala 16:16]
  reg [255:0] mem_7; // @[Ram.scala 16:16]
  reg [255:0] mem_8; // @[Ram.scala 16:16]
  reg [255:0] mem_9; // @[Ram.scala 16:16]
  reg [255:0] mem_10; // @[Ram.scala 16:16]
  reg [255:0] mem_11; // @[Ram.scala 16:16]
  reg [255:0] mem_12; // @[Ram.scala 16:16]
  reg [255:0] mem_13; // @[Ram.scala 16:16]
  reg [255:0] mem_14; // @[Ram.scala 16:16]
  reg [255:0] mem_15; // @[Ram.scala 16:16]
  reg [255:0] mem_16; // @[Ram.scala 16:16]
  reg [255:0] mem_17; // @[Ram.scala 16:16]
  reg [255:0] mem_18; // @[Ram.scala 16:16]
  reg [255:0] mem_19; // @[Ram.scala 16:16]
  reg [255:0] mem_20; // @[Ram.scala 16:16]
  reg [255:0] mem_21; // @[Ram.scala 16:16]
  reg [255:0] mem_22; // @[Ram.scala 16:16]
  reg [255:0] mem_23; // @[Ram.scala 16:16]
  reg [255:0] mem_24; // @[Ram.scala 16:16]
  reg [255:0] mem_25; // @[Ram.scala 16:16]
  reg [255:0] mem_26; // @[Ram.scala 16:16]
  reg [255:0] mem_27; // @[Ram.scala 16:16]
  reg [255:0] mem_28; // @[Ram.scala 16:16]
  reg [255:0] mem_29; // @[Ram.scala 16:16]
  reg [255:0] mem_30; // @[Ram.scala 16:16]
  reg [255:0] mem_31; // @[Ram.scala 16:16]
  reg [255:0] mem_32; // @[Ram.scala 16:16]
  reg [255:0] mem_33; // @[Ram.scala 16:16]
  reg [255:0] mem_34; // @[Ram.scala 16:16]
  reg [255:0] mem_35; // @[Ram.scala 16:16]
  reg [255:0] mem_36; // @[Ram.scala 16:16]
  reg [255:0] mem_37; // @[Ram.scala 16:16]
  reg [255:0] mem_38; // @[Ram.scala 16:16]
  reg [255:0] mem_39; // @[Ram.scala 16:16]
  reg [255:0] mem_40; // @[Ram.scala 16:16]
  reg [255:0] mem_41; // @[Ram.scala 16:16]
  reg [255:0] mem_42; // @[Ram.scala 16:16]
  reg [255:0] mem_43; // @[Ram.scala 16:16]
  reg [255:0] mem_44; // @[Ram.scala 16:16]
  reg [255:0] mem_45; // @[Ram.scala 16:16]
  reg [255:0] mem_46; // @[Ram.scala 16:16]
  reg [255:0] mem_47; // @[Ram.scala 16:16]
  reg [255:0] mem_48; // @[Ram.scala 16:16]
  reg [255:0] mem_49; // @[Ram.scala 16:16]
  reg [255:0] mem_50; // @[Ram.scala 16:16]
  reg [255:0] mem_51; // @[Ram.scala 16:16]
  reg [255:0] mem_52; // @[Ram.scala 16:16]
  reg [255:0] mem_53; // @[Ram.scala 16:16]
  reg [255:0] mem_54; // @[Ram.scala 16:16]
  reg [255:0] mem_55; // @[Ram.scala 16:16]
  reg [255:0] mem_56; // @[Ram.scala 16:16]
  reg [255:0] mem_57; // @[Ram.scala 16:16]
  reg [255:0] mem_58; // @[Ram.scala 16:16]
  reg [255:0] mem_59; // @[Ram.scala 16:16]
  reg [255:0] mem_60; // @[Ram.scala 16:16]
  reg [255:0] mem_61; // @[Ram.scala 16:16]
  reg [255:0] mem_62; // @[Ram.scala 16:16]
  reg [255:0] mem_63; // @[Ram.scala 16:16]
  reg [255:0] mem_64; // @[Ram.scala 16:16]
  reg [255:0] mem_65; // @[Ram.scala 16:16]
  reg [255:0] mem_66; // @[Ram.scala 16:16]
  reg [255:0] mem_67; // @[Ram.scala 16:16]
  reg [255:0] mem_68; // @[Ram.scala 16:16]
  reg [255:0] mem_69; // @[Ram.scala 16:16]
  reg [255:0] mem_70; // @[Ram.scala 16:16]
  reg [255:0] mem_71; // @[Ram.scala 16:16]
  reg [255:0] mem_72; // @[Ram.scala 16:16]
  reg [255:0] mem_73; // @[Ram.scala 16:16]
  reg [255:0] mem_74; // @[Ram.scala 16:16]
  reg [255:0] mem_75; // @[Ram.scala 16:16]
  reg [255:0] mem_76; // @[Ram.scala 16:16]
  reg [255:0] mem_77; // @[Ram.scala 16:16]
  reg [255:0] mem_78; // @[Ram.scala 16:16]
  reg [255:0] mem_79; // @[Ram.scala 16:16]
  reg [255:0] mem_80; // @[Ram.scala 16:16]
  reg [255:0] mem_81; // @[Ram.scala 16:16]
  reg [255:0] mem_82; // @[Ram.scala 16:16]
  reg [255:0] mem_83; // @[Ram.scala 16:16]
  reg [255:0] mem_84; // @[Ram.scala 16:16]
  reg [255:0] mem_85; // @[Ram.scala 16:16]
  reg [255:0] mem_86; // @[Ram.scala 16:16]
  reg [255:0] mem_87; // @[Ram.scala 16:16]
  reg [255:0] mem_88; // @[Ram.scala 16:16]
  reg [255:0] mem_89; // @[Ram.scala 16:16]
  reg [255:0] mem_90; // @[Ram.scala 16:16]
  reg [255:0] mem_91; // @[Ram.scala 16:16]
  reg [255:0] mem_92; // @[Ram.scala 16:16]
  reg [255:0] mem_93; // @[Ram.scala 16:16]
  reg [255:0] mem_94; // @[Ram.scala 16:16]
  reg [255:0] mem_95; // @[Ram.scala 16:16]
  reg [255:0] mem_96; // @[Ram.scala 16:16]
  reg [255:0] mem_97; // @[Ram.scala 16:16]
  reg [255:0] mem_98; // @[Ram.scala 16:16]
  reg [255:0] mem_99; // @[Ram.scala 16:16]
  reg [255:0] mem_100; // @[Ram.scala 16:16]
  reg [255:0] mem_101; // @[Ram.scala 16:16]
  reg [255:0] mem_102; // @[Ram.scala 16:16]
  reg [255:0] mem_103; // @[Ram.scala 16:16]
  reg [255:0] mem_104; // @[Ram.scala 16:16]
  reg [255:0] mem_105; // @[Ram.scala 16:16]
  reg [255:0] mem_106; // @[Ram.scala 16:16]
  reg [255:0] mem_107; // @[Ram.scala 16:16]
  reg [255:0] mem_108; // @[Ram.scala 16:16]
  reg [255:0] mem_109; // @[Ram.scala 16:16]
  reg [255:0] mem_110; // @[Ram.scala 16:16]
  reg [255:0] mem_111; // @[Ram.scala 16:16]
  reg [255:0] mem_112; // @[Ram.scala 16:16]
  reg [255:0] mem_113; // @[Ram.scala 16:16]
  reg [255:0] mem_114; // @[Ram.scala 16:16]
  reg [255:0] mem_115; // @[Ram.scala 16:16]
  reg [255:0] mem_116; // @[Ram.scala 16:16]
  reg [255:0] mem_117; // @[Ram.scala 16:16]
  reg [255:0] mem_118; // @[Ram.scala 16:16]
  reg [255:0] mem_119; // @[Ram.scala 16:16]
  reg [255:0] mem_120; // @[Ram.scala 16:16]
  reg [255:0] mem_121; // @[Ram.scala 16:16]
  reg [255:0] mem_122; // @[Ram.scala 16:16]
  reg [255:0] mem_123; // @[Ram.scala 16:16]
  reg [255:0] mem_124; // @[Ram.scala 16:16]
  reg [255:0] mem_125; // @[Ram.scala 16:16]
  reg [255:0] mem_126; // @[Ram.scala 16:16]
  reg [255:0] mem_127; // @[Ram.scala 16:16]
  reg [255:0] mem_128; // @[Ram.scala 16:16]
  reg [255:0] mem_129; // @[Ram.scala 16:16]
  reg [255:0] mem_130; // @[Ram.scala 16:16]
  reg [255:0] mem_131; // @[Ram.scala 16:16]
  reg [255:0] mem_132; // @[Ram.scala 16:16]
  reg [255:0] mem_133; // @[Ram.scala 16:16]
  reg [255:0] mem_134; // @[Ram.scala 16:16]
  reg [255:0] mem_135; // @[Ram.scala 16:16]
  reg [255:0] mem_136; // @[Ram.scala 16:16]
  reg [255:0] mem_137; // @[Ram.scala 16:16]
  reg [255:0] mem_138; // @[Ram.scala 16:16]
  reg [255:0] mem_139; // @[Ram.scala 16:16]
  reg [255:0] mem_140; // @[Ram.scala 16:16]
  reg [255:0] mem_141; // @[Ram.scala 16:16]
  reg [255:0] mem_142; // @[Ram.scala 16:16]
  reg [255:0] mem_143; // @[Ram.scala 16:16]
  reg [255:0] mem_144; // @[Ram.scala 16:16]
  reg [255:0] mem_145; // @[Ram.scala 16:16]
  reg [255:0] mem_146; // @[Ram.scala 16:16]
  reg [255:0] mem_147; // @[Ram.scala 16:16]
  reg [255:0] mem_148; // @[Ram.scala 16:16]
  reg [255:0] mem_149; // @[Ram.scala 16:16]
  reg [255:0] mem_150; // @[Ram.scala 16:16]
  reg [255:0] mem_151; // @[Ram.scala 16:16]
  reg [255:0] mem_152; // @[Ram.scala 16:16]
  reg [255:0] mem_153; // @[Ram.scala 16:16]
  reg [255:0] mem_154; // @[Ram.scala 16:16]
  reg [255:0] mem_155; // @[Ram.scala 16:16]
  reg [255:0] mem_156; // @[Ram.scala 16:16]
  reg [255:0] mem_157; // @[Ram.scala 16:16]
  reg [255:0] mem_158; // @[Ram.scala 16:16]
  reg [255:0] mem_159; // @[Ram.scala 16:16]
  reg [255:0] mem_160; // @[Ram.scala 16:16]
  reg [255:0] mem_161; // @[Ram.scala 16:16]
  reg [255:0] mem_162; // @[Ram.scala 16:16]
  reg [255:0] mem_163; // @[Ram.scala 16:16]
  reg [255:0] mem_164; // @[Ram.scala 16:16]
  reg [255:0] mem_165; // @[Ram.scala 16:16]
  reg [255:0] mem_166; // @[Ram.scala 16:16]
  reg [255:0] mem_167; // @[Ram.scala 16:16]
  reg [255:0] mem_168; // @[Ram.scala 16:16]
  reg [255:0] mem_169; // @[Ram.scala 16:16]
  reg [255:0] mem_170; // @[Ram.scala 16:16]
  reg [255:0] mem_171; // @[Ram.scala 16:16]
  reg [255:0] mem_172; // @[Ram.scala 16:16]
  reg [255:0] mem_173; // @[Ram.scala 16:16]
  reg [255:0] mem_174; // @[Ram.scala 16:16]
  reg [255:0] mem_175; // @[Ram.scala 16:16]
  reg [255:0] mem_176; // @[Ram.scala 16:16]
  reg [255:0] mem_177; // @[Ram.scala 16:16]
  reg [255:0] mem_178; // @[Ram.scala 16:16]
  reg [255:0] mem_179; // @[Ram.scala 16:16]
  reg [255:0] mem_180; // @[Ram.scala 16:16]
  reg [255:0] mem_181; // @[Ram.scala 16:16]
  reg [255:0] mem_182; // @[Ram.scala 16:16]
  reg [255:0] mem_183; // @[Ram.scala 16:16]
  reg [255:0] mem_184; // @[Ram.scala 16:16]
  reg [255:0] mem_185; // @[Ram.scala 16:16]
  reg [255:0] mem_186; // @[Ram.scala 16:16]
  reg [255:0] mem_187; // @[Ram.scala 16:16]
  reg [255:0] mem_188; // @[Ram.scala 16:16]
  reg [255:0] mem_189; // @[Ram.scala 16:16]
  reg [255:0] mem_190; // @[Ram.scala 16:16]
  reg [255:0] mem_191; // @[Ram.scala 16:16]
  reg [255:0] mem_192; // @[Ram.scala 16:16]
  reg [255:0] mem_193; // @[Ram.scala 16:16]
  reg [255:0] mem_194; // @[Ram.scala 16:16]
  reg [255:0] mem_195; // @[Ram.scala 16:16]
  reg [255:0] mem_196; // @[Ram.scala 16:16]
  reg [255:0] mem_197; // @[Ram.scala 16:16]
  reg [255:0] mem_198; // @[Ram.scala 16:16]
  reg [255:0] mem_199; // @[Ram.scala 16:16]
  reg [255:0] mem_200; // @[Ram.scala 16:16]
  reg [255:0] mem_201; // @[Ram.scala 16:16]
  reg [255:0] mem_202; // @[Ram.scala 16:16]
  reg [255:0] mem_203; // @[Ram.scala 16:16]
  reg [255:0] mem_204; // @[Ram.scala 16:16]
  reg [255:0] mem_205; // @[Ram.scala 16:16]
  reg [255:0] mem_206; // @[Ram.scala 16:16]
  reg [255:0] mem_207; // @[Ram.scala 16:16]
  reg [255:0] mem_208; // @[Ram.scala 16:16]
  reg [255:0] mem_209; // @[Ram.scala 16:16]
  reg [255:0] mem_210; // @[Ram.scala 16:16]
  reg [255:0] mem_211; // @[Ram.scala 16:16]
  reg [255:0] mem_212; // @[Ram.scala 16:16]
  reg [255:0] mem_213; // @[Ram.scala 16:16]
  reg [255:0] mem_214; // @[Ram.scala 16:16]
  reg [255:0] mem_215; // @[Ram.scala 16:16]
  reg [255:0] mem_216; // @[Ram.scala 16:16]
  reg [255:0] mem_217; // @[Ram.scala 16:16]
  reg [255:0] mem_218; // @[Ram.scala 16:16]
  reg [255:0] mem_219; // @[Ram.scala 16:16]
  reg [255:0] mem_220; // @[Ram.scala 16:16]
  reg [255:0] mem_221; // @[Ram.scala 16:16]
  reg [255:0] mem_222; // @[Ram.scala 16:16]
  reg [255:0] mem_223; // @[Ram.scala 16:16]
  reg [255:0] mem_224; // @[Ram.scala 16:16]
  reg [255:0] mem_225; // @[Ram.scala 16:16]
  reg [255:0] mem_226; // @[Ram.scala 16:16]
  reg [255:0] mem_227; // @[Ram.scala 16:16]
  reg [255:0] mem_228; // @[Ram.scala 16:16]
  reg [255:0] mem_229; // @[Ram.scala 16:16]
  reg [255:0] mem_230; // @[Ram.scala 16:16]
  reg [255:0] mem_231; // @[Ram.scala 16:16]
  reg [255:0] mem_232; // @[Ram.scala 16:16]
  reg [255:0] mem_233; // @[Ram.scala 16:16]
  reg [255:0] mem_234; // @[Ram.scala 16:16]
  reg [255:0] mem_235; // @[Ram.scala 16:16]
  reg [255:0] mem_236; // @[Ram.scala 16:16]
  reg [255:0] mem_237; // @[Ram.scala 16:16]
  reg [255:0] mem_238; // @[Ram.scala 16:16]
  reg [255:0] mem_239; // @[Ram.scala 16:16]
  reg [255:0] mem_240; // @[Ram.scala 16:16]
  reg [255:0] mem_241; // @[Ram.scala 16:16]
  reg [255:0] mem_242; // @[Ram.scala 16:16]
  reg [255:0] mem_243; // @[Ram.scala 16:16]
  reg [255:0] mem_244; // @[Ram.scala 16:16]
  reg [255:0] mem_245; // @[Ram.scala 16:16]
  reg [255:0] mem_246; // @[Ram.scala 16:16]
  reg [255:0] mem_247; // @[Ram.scala 16:16]
  reg [255:0] mem_248; // @[Ram.scala 16:16]
  reg [255:0] mem_249; // @[Ram.scala 16:16]
  reg [255:0] mem_250; // @[Ram.scala 16:16]
  reg [255:0] mem_251; // @[Ram.scala 16:16]
  reg [255:0] mem_252; // @[Ram.scala 16:16]
  reg [255:0] mem_253; // @[Ram.scala 16:16]
  reg [255:0] mem_254; // @[Ram.scala 16:16]
  reg [255:0] mem_255; // @[Ram.scala 16:16]
  reg [255:0] mem_256; // @[Ram.scala 16:16]
  reg [255:0] mem_257; // @[Ram.scala 16:16]
  reg [255:0] mem_258; // @[Ram.scala 16:16]
  reg [255:0] mem_259; // @[Ram.scala 16:16]
  reg [255:0] mem_260; // @[Ram.scala 16:16]
  reg [255:0] mem_261; // @[Ram.scala 16:16]
  reg [255:0] mem_262; // @[Ram.scala 16:16]
  reg [255:0] mem_263; // @[Ram.scala 16:16]
  reg [255:0] mem_264; // @[Ram.scala 16:16]
  reg [255:0] mem_265; // @[Ram.scala 16:16]
  reg [255:0] mem_266; // @[Ram.scala 16:16]
  reg [255:0] mem_267; // @[Ram.scala 16:16]
  reg [255:0] mem_268; // @[Ram.scala 16:16]
  reg [255:0] mem_269; // @[Ram.scala 16:16]
  reg [255:0] mem_270; // @[Ram.scala 16:16]
  reg [255:0] mem_271; // @[Ram.scala 16:16]
  reg [255:0] mem_272; // @[Ram.scala 16:16]
  reg [255:0] mem_273; // @[Ram.scala 16:16]
  reg [255:0] mem_274; // @[Ram.scala 16:16]
  reg [255:0] mem_275; // @[Ram.scala 16:16]
  reg [255:0] mem_276; // @[Ram.scala 16:16]
  reg [255:0] mem_277; // @[Ram.scala 16:16]
  reg [255:0] mem_278; // @[Ram.scala 16:16]
  reg [255:0] mem_279; // @[Ram.scala 16:16]
  reg [255:0] mem_280; // @[Ram.scala 16:16]
  reg [255:0] mem_281; // @[Ram.scala 16:16]
  reg [255:0] mem_282; // @[Ram.scala 16:16]
  reg [255:0] mem_283; // @[Ram.scala 16:16]
  reg [255:0] mem_284; // @[Ram.scala 16:16]
  reg [255:0] mem_285; // @[Ram.scala 16:16]
  reg [255:0] mem_286; // @[Ram.scala 16:16]
  reg [255:0] mem_287; // @[Ram.scala 16:16]
  reg [255:0] mem_288; // @[Ram.scala 16:16]
  reg [255:0] mem_289; // @[Ram.scala 16:16]
  reg [255:0] mem_290; // @[Ram.scala 16:16]
  reg [255:0] mem_291; // @[Ram.scala 16:16]
  reg [255:0] mem_292; // @[Ram.scala 16:16]
  reg [255:0] mem_293; // @[Ram.scala 16:16]
  reg [255:0] mem_294; // @[Ram.scala 16:16]
  reg [255:0] mem_295; // @[Ram.scala 16:16]
  reg [255:0] mem_296; // @[Ram.scala 16:16]
  reg [255:0] mem_297; // @[Ram.scala 16:16]
  reg [255:0] mem_298; // @[Ram.scala 16:16]
  reg [255:0] mem_299; // @[Ram.scala 16:16]
  reg [255:0] mem_300; // @[Ram.scala 16:16]
  reg [255:0] mem_301; // @[Ram.scala 16:16]
  reg [255:0] mem_302; // @[Ram.scala 16:16]
  reg [255:0] mem_303; // @[Ram.scala 16:16]
  reg [255:0] mem_304; // @[Ram.scala 16:16]
  reg [255:0] mem_305; // @[Ram.scala 16:16]
  reg [255:0] mem_306; // @[Ram.scala 16:16]
  reg [255:0] mem_307; // @[Ram.scala 16:16]
  reg [255:0] mem_308; // @[Ram.scala 16:16]
  reg [255:0] mem_309; // @[Ram.scala 16:16]
  reg [255:0] mem_310; // @[Ram.scala 16:16]
  reg [255:0] mem_311; // @[Ram.scala 16:16]
  reg [255:0] mem_312; // @[Ram.scala 16:16]
  reg [255:0] mem_313; // @[Ram.scala 16:16]
  reg [255:0] mem_314; // @[Ram.scala 16:16]
  reg [255:0] mem_315; // @[Ram.scala 16:16]
  reg [255:0] mem_316; // @[Ram.scala 16:16]
  reg [255:0] mem_317; // @[Ram.scala 16:16]
  reg [255:0] mem_318; // @[Ram.scala 16:16]
  reg [255:0] mem_319; // @[Ram.scala 16:16]
  reg [255:0] mem_320; // @[Ram.scala 16:16]
  reg [255:0] mem_321; // @[Ram.scala 16:16]
  reg [255:0] mem_322; // @[Ram.scala 16:16]
  reg [255:0] mem_323; // @[Ram.scala 16:16]
  reg [255:0] mem_324; // @[Ram.scala 16:16]
  reg [255:0] mem_325; // @[Ram.scala 16:16]
  reg [255:0] mem_326; // @[Ram.scala 16:16]
  reg [255:0] mem_327; // @[Ram.scala 16:16]
  reg [255:0] mem_328; // @[Ram.scala 16:16]
  reg [255:0] mem_329; // @[Ram.scala 16:16]
  reg [255:0] mem_330; // @[Ram.scala 16:16]
  reg [255:0] mem_331; // @[Ram.scala 16:16]
  reg [255:0] mem_332; // @[Ram.scala 16:16]
  reg [255:0] mem_333; // @[Ram.scala 16:16]
  reg [255:0] mem_334; // @[Ram.scala 16:16]
  reg [255:0] mem_335; // @[Ram.scala 16:16]
  reg [255:0] mem_336; // @[Ram.scala 16:16]
  reg [255:0] mem_337; // @[Ram.scala 16:16]
  reg [255:0] mem_338; // @[Ram.scala 16:16]
  reg [255:0] mem_339; // @[Ram.scala 16:16]
  reg [255:0] mem_340; // @[Ram.scala 16:16]
  reg [255:0] mem_341; // @[Ram.scala 16:16]
  reg [255:0] mem_342; // @[Ram.scala 16:16]
  reg [255:0] mem_343; // @[Ram.scala 16:16]
  reg [255:0] mem_344; // @[Ram.scala 16:16]
  reg [255:0] mem_345; // @[Ram.scala 16:16]
  reg [255:0] mem_346; // @[Ram.scala 16:16]
  reg [255:0] mem_347; // @[Ram.scala 16:16]
  reg [255:0] mem_348; // @[Ram.scala 16:16]
  reg [255:0] mem_349; // @[Ram.scala 16:16]
  reg [255:0] mem_350; // @[Ram.scala 16:16]
  reg [255:0] mem_351; // @[Ram.scala 16:16]
  reg [255:0] mem_352; // @[Ram.scala 16:16]
  reg [255:0] mem_353; // @[Ram.scala 16:16]
  reg [255:0] mem_354; // @[Ram.scala 16:16]
  reg [255:0] mem_355; // @[Ram.scala 16:16]
  reg [255:0] mem_356; // @[Ram.scala 16:16]
  reg [255:0] mem_357; // @[Ram.scala 16:16]
  reg [255:0] mem_358; // @[Ram.scala 16:16]
  reg [255:0] mem_359; // @[Ram.scala 16:16]
  reg [255:0] mem_360; // @[Ram.scala 16:16]
  reg [255:0] mem_361; // @[Ram.scala 16:16]
  reg [255:0] mem_362; // @[Ram.scala 16:16]
  reg [255:0] mem_363; // @[Ram.scala 16:16]
  reg [255:0] mem_364; // @[Ram.scala 16:16]
  reg [255:0] mem_365; // @[Ram.scala 16:16]
  reg [255:0] mem_366; // @[Ram.scala 16:16]
  reg [255:0] mem_367; // @[Ram.scala 16:16]
  reg [255:0] mem_368; // @[Ram.scala 16:16]
  reg [255:0] mem_369; // @[Ram.scala 16:16]
  reg [255:0] mem_370; // @[Ram.scala 16:16]
  reg [255:0] mem_371; // @[Ram.scala 16:16]
  reg [255:0] mem_372; // @[Ram.scala 16:16]
  reg [255:0] mem_373; // @[Ram.scala 16:16]
  reg [255:0] mem_374; // @[Ram.scala 16:16]
  reg [255:0] mem_375; // @[Ram.scala 16:16]
  reg [255:0] mem_376; // @[Ram.scala 16:16]
  reg [255:0] mem_377; // @[Ram.scala 16:16]
  reg [255:0] mem_378; // @[Ram.scala 16:16]
  reg [255:0] mem_379; // @[Ram.scala 16:16]
  reg [255:0] mem_380; // @[Ram.scala 16:16]
  reg [255:0] mem_381; // @[Ram.scala 16:16]
  reg [255:0] mem_382; // @[Ram.scala 16:16]
  reg [255:0] mem_383; // @[Ram.scala 16:16]
  reg [255:0] mem_384; // @[Ram.scala 16:16]
  reg [255:0] mem_385; // @[Ram.scala 16:16]
  reg [255:0] mem_386; // @[Ram.scala 16:16]
  reg [255:0] mem_387; // @[Ram.scala 16:16]
  reg [255:0] mem_388; // @[Ram.scala 16:16]
  reg [255:0] mem_389; // @[Ram.scala 16:16]
  reg [255:0] mem_390; // @[Ram.scala 16:16]
  reg [255:0] mem_391; // @[Ram.scala 16:16]
  reg [255:0] mem_392; // @[Ram.scala 16:16]
  reg [255:0] mem_393; // @[Ram.scala 16:16]
  reg [255:0] mem_394; // @[Ram.scala 16:16]
  reg [255:0] mem_395; // @[Ram.scala 16:16]
  reg [255:0] mem_396; // @[Ram.scala 16:16]
  reg [255:0] mem_397; // @[Ram.scala 16:16]
  reg [255:0] mem_398; // @[Ram.scala 16:16]
  reg [255:0] mem_399; // @[Ram.scala 16:16]
  reg [255:0] mem_400; // @[Ram.scala 16:16]
  reg [255:0] mem_401; // @[Ram.scala 16:16]
  reg [255:0] mem_402; // @[Ram.scala 16:16]
  reg [255:0] mem_403; // @[Ram.scala 16:16]
  reg [255:0] mem_404; // @[Ram.scala 16:16]
  reg [255:0] mem_405; // @[Ram.scala 16:16]
  reg [255:0] mem_406; // @[Ram.scala 16:16]
  reg [255:0] mem_407; // @[Ram.scala 16:16]
  reg [255:0] mem_408; // @[Ram.scala 16:16]
  reg [255:0] mem_409; // @[Ram.scala 16:16]
  reg [255:0] mem_410; // @[Ram.scala 16:16]
  reg [255:0] mem_411; // @[Ram.scala 16:16]
  reg [255:0] mem_412; // @[Ram.scala 16:16]
  reg [255:0] mem_413; // @[Ram.scala 16:16]
  reg [255:0] mem_414; // @[Ram.scala 16:16]
  reg [255:0] mem_415; // @[Ram.scala 16:16]
  reg [255:0] mem_416; // @[Ram.scala 16:16]
  reg [255:0] mem_417; // @[Ram.scala 16:16]
  reg [255:0] mem_418; // @[Ram.scala 16:16]
  reg [255:0] mem_419; // @[Ram.scala 16:16]
  reg [255:0] mem_420; // @[Ram.scala 16:16]
  reg [255:0] mem_421; // @[Ram.scala 16:16]
  reg [255:0] mem_422; // @[Ram.scala 16:16]
  reg [255:0] mem_423; // @[Ram.scala 16:16]
  reg [255:0] mem_424; // @[Ram.scala 16:16]
  reg [255:0] mem_425; // @[Ram.scala 16:16]
  reg [255:0] mem_426; // @[Ram.scala 16:16]
  reg [255:0] mem_427; // @[Ram.scala 16:16]
  reg [255:0] mem_428; // @[Ram.scala 16:16]
  reg [255:0] mem_429; // @[Ram.scala 16:16]
  reg [255:0] mem_430; // @[Ram.scala 16:16]
  reg [255:0] mem_431; // @[Ram.scala 16:16]
  reg [255:0] mem_432; // @[Ram.scala 16:16]
  reg [255:0] mem_433; // @[Ram.scala 16:16]
  reg [255:0] mem_434; // @[Ram.scala 16:16]
  reg [255:0] mem_435; // @[Ram.scala 16:16]
  reg [255:0] mem_436; // @[Ram.scala 16:16]
  reg [255:0] mem_437; // @[Ram.scala 16:16]
  reg [255:0] mem_438; // @[Ram.scala 16:16]
  reg [255:0] mem_439; // @[Ram.scala 16:16]
  reg [255:0] mem_440; // @[Ram.scala 16:16]
  reg [255:0] mem_441; // @[Ram.scala 16:16]
  reg [255:0] mem_442; // @[Ram.scala 16:16]
  reg [255:0] mem_443; // @[Ram.scala 16:16]
  reg [255:0] mem_444; // @[Ram.scala 16:16]
  reg [255:0] mem_445; // @[Ram.scala 16:16]
  reg [255:0] mem_446; // @[Ram.scala 16:16]
  reg [255:0] mem_447; // @[Ram.scala 16:16]
  reg [255:0] mem_448; // @[Ram.scala 16:16]
  reg [255:0] mem_449; // @[Ram.scala 16:16]
  reg [255:0] mem_450; // @[Ram.scala 16:16]
  reg [255:0] mem_451; // @[Ram.scala 16:16]
  reg [255:0] mem_452; // @[Ram.scala 16:16]
  reg [255:0] mem_453; // @[Ram.scala 16:16]
  reg [255:0] mem_454; // @[Ram.scala 16:16]
  reg [255:0] mem_455; // @[Ram.scala 16:16]
  reg [255:0] mem_456; // @[Ram.scala 16:16]
  reg [255:0] mem_457; // @[Ram.scala 16:16]
  reg [255:0] mem_458; // @[Ram.scala 16:16]
  reg [255:0] mem_459; // @[Ram.scala 16:16]
  reg [255:0] mem_460; // @[Ram.scala 16:16]
  reg [255:0] mem_461; // @[Ram.scala 16:16]
  reg [255:0] mem_462; // @[Ram.scala 16:16]
  reg [255:0] mem_463; // @[Ram.scala 16:16]
  reg [255:0] mem_464; // @[Ram.scala 16:16]
  reg [255:0] mem_465; // @[Ram.scala 16:16]
  reg [255:0] mem_466; // @[Ram.scala 16:16]
  reg [255:0] mem_467; // @[Ram.scala 16:16]
  reg [255:0] mem_468; // @[Ram.scala 16:16]
  reg [255:0] mem_469; // @[Ram.scala 16:16]
  reg [255:0] mem_470; // @[Ram.scala 16:16]
  reg [255:0] mem_471; // @[Ram.scala 16:16]
  reg [255:0] mem_472; // @[Ram.scala 16:16]
  reg [255:0] mem_473; // @[Ram.scala 16:16]
  reg [255:0] mem_474; // @[Ram.scala 16:16]
  reg [255:0] mem_475; // @[Ram.scala 16:16]
  reg [255:0] mem_476; // @[Ram.scala 16:16]
  reg [255:0] mem_477; // @[Ram.scala 16:16]
  reg [255:0] mem_478; // @[Ram.scala 16:16]
  reg [255:0] mem_479; // @[Ram.scala 16:16]
  reg [255:0] mem_480; // @[Ram.scala 16:16]
  reg [255:0] mem_481; // @[Ram.scala 16:16]
  reg [255:0] mem_482; // @[Ram.scala 16:16]
  reg [255:0] mem_483; // @[Ram.scala 16:16]
  reg [255:0] mem_484; // @[Ram.scala 16:16]
  reg [255:0] mem_485; // @[Ram.scala 16:16]
  reg [255:0] mem_486; // @[Ram.scala 16:16]
  reg [255:0] mem_487; // @[Ram.scala 16:16]
  reg [255:0] mem_488; // @[Ram.scala 16:16]
  reg [255:0] mem_489; // @[Ram.scala 16:16]
  reg [255:0] mem_490; // @[Ram.scala 16:16]
  reg [255:0] mem_491; // @[Ram.scala 16:16]
  reg [255:0] mem_492; // @[Ram.scala 16:16]
  reg [255:0] mem_493; // @[Ram.scala 16:16]
  reg [255:0] mem_494; // @[Ram.scala 16:16]
  reg [255:0] mem_495; // @[Ram.scala 16:16]
  reg [255:0] mem_496; // @[Ram.scala 16:16]
  reg [255:0] mem_497; // @[Ram.scala 16:16]
  reg [255:0] mem_498; // @[Ram.scala 16:16]
  reg [255:0] mem_499; // @[Ram.scala 16:16]
  reg [255:0] mem_500; // @[Ram.scala 16:16]
  reg [255:0] mem_501; // @[Ram.scala 16:16]
  reg [255:0] mem_502; // @[Ram.scala 16:16]
  reg [255:0] mem_503; // @[Ram.scala 16:16]
  reg [255:0] mem_504; // @[Ram.scala 16:16]
  reg [255:0] mem_505; // @[Ram.scala 16:16]
  reg [255:0] mem_506; // @[Ram.scala 16:16]
  reg [255:0] mem_507; // @[Ram.scala 16:16]
  reg [255:0] mem_508; // @[Ram.scala 16:16]
  reg [255:0] mem_509; // @[Ram.scala 16:16]
  reg [255:0] mem_510; // @[Ram.scala 16:16]
  reg [255:0] mem_511; // @[Ram.scala 16:16]
  reg [255:0] mem_512; // @[Ram.scala 16:16]
  reg [255:0] mem_513; // @[Ram.scala 16:16]
  reg [255:0] mem_514; // @[Ram.scala 16:16]
  reg [255:0] mem_515; // @[Ram.scala 16:16]
  reg [255:0] mem_516; // @[Ram.scala 16:16]
  reg [255:0] mem_517; // @[Ram.scala 16:16]
  reg [255:0] mem_518; // @[Ram.scala 16:16]
  reg [255:0] mem_519; // @[Ram.scala 16:16]
  reg [255:0] mem_520; // @[Ram.scala 16:16]
  reg [255:0] mem_521; // @[Ram.scala 16:16]
  reg [255:0] mem_522; // @[Ram.scala 16:16]
  reg [255:0] mem_523; // @[Ram.scala 16:16]
  reg [255:0] mem_524; // @[Ram.scala 16:16]
  reg [255:0] mem_525; // @[Ram.scala 16:16]
  reg [255:0] mem_526; // @[Ram.scala 16:16]
  reg [255:0] mem_527; // @[Ram.scala 16:16]
  reg [255:0] mem_528; // @[Ram.scala 16:16]
  reg [255:0] mem_529; // @[Ram.scala 16:16]
  reg [255:0] mem_530; // @[Ram.scala 16:16]
  reg [255:0] mem_531; // @[Ram.scala 16:16]
  reg [255:0] mem_532; // @[Ram.scala 16:16]
  reg [255:0] mem_533; // @[Ram.scala 16:16]
  reg [255:0] mem_534; // @[Ram.scala 16:16]
  reg [255:0] mem_535; // @[Ram.scala 16:16]
  reg [255:0] mem_536; // @[Ram.scala 16:16]
  reg [255:0] mem_537; // @[Ram.scala 16:16]
  reg [255:0] mem_538; // @[Ram.scala 16:16]
  reg [255:0] mem_539; // @[Ram.scala 16:16]
  reg [255:0] mem_540; // @[Ram.scala 16:16]
  reg [255:0] mem_541; // @[Ram.scala 16:16]
  reg [255:0] mem_542; // @[Ram.scala 16:16]
  reg [255:0] mem_543; // @[Ram.scala 16:16]
  reg [255:0] mem_544; // @[Ram.scala 16:16]
  reg [255:0] mem_545; // @[Ram.scala 16:16]
  reg [255:0] mem_546; // @[Ram.scala 16:16]
  reg [255:0] mem_547; // @[Ram.scala 16:16]
  reg [255:0] mem_548; // @[Ram.scala 16:16]
  reg [255:0] mem_549; // @[Ram.scala 16:16]
  reg [255:0] mem_550; // @[Ram.scala 16:16]
  reg [255:0] mem_551; // @[Ram.scala 16:16]
  reg [255:0] mem_552; // @[Ram.scala 16:16]
  reg [255:0] mem_553; // @[Ram.scala 16:16]
  reg [255:0] mem_554; // @[Ram.scala 16:16]
  reg [255:0] mem_555; // @[Ram.scala 16:16]
  reg [255:0] mem_556; // @[Ram.scala 16:16]
  reg [255:0] mem_557; // @[Ram.scala 16:16]
  reg [255:0] mem_558; // @[Ram.scala 16:16]
  reg [255:0] mem_559; // @[Ram.scala 16:16]
  reg [255:0] mem_560; // @[Ram.scala 16:16]
  reg [255:0] mem_561; // @[Ram.scala 16:16]
  reg [255:0] mem_562; // @[Ram.scala 16:16]
  reg [255:0] mem_563; // @[Ram.scala 16:16]
  reg [255:0] mem_564; // @[Ram.scala 16:16]
  reg [255:0] mem_565; // @[Ram.scala 16:16]
  reg [255:0] mem_566; // @[Ram.scala 16:16]
  reg [255:0] mem_567; // @[Ram.scala 16:16]
  reg [255:0] mem_568; // @[Ram.scala 16:16]
  reg [255:0] mem_569; // @[Ram.scala 16:16]
  reg [255:0] mem_570; // @[Ram.scala 16:16]
  reg [255:0] mem_571; // @[Ram.scala 16:16]
  reg [255:0] mem_572; // @[Ram.scala 16:16]
  reg [255:0] mem_573; // @[Ram.scala 16:16]
  reg [255:0] mem_574; // @[Ram.scala 16:16]
  reg [255:0] mem_575; // @[Ram.scala 16:16]
  reg [255:0] mem_576; // @[Ram.scala 16:16]
  reg [255:0] mem_577; // @[Ram.scala 16:16]
  reg [255:0] mem_578; // @[Ram.scala 16:16]
  reg [255:0] mem_579; // @[Ram.scala 16:16]
  reg [255:0] mem_580; // @[Ram.scala 16:16]
  reg [255:0] mem_581; // @[Ram.scala 16:16]
  reg [255:0] mem_582; // @[Ram.scala 16:16]
  reg [255:0] mem_583; // @[Ram.scala 16:16]
  reg [255:0] mem_584; // @[Ram.scala 16:16]
  reg [255:0] mem_585; // @[Ram.scala 16:16]
  reg [255:0] mem_586; // @[Ram.scala 16:16]
  reg [255:0] mem_587; // @[Ram.scala 16:16]
  reg [255:0] mem_588; // @[Ram.scala 16:16]
  reg [255:0] mem_589; // @[Ram.scala 16:16]
  reg [255:0] mem_590; // @[Ram.scala 16:16]
  reg [255:0] mem_591; // @[Ram.scala 16:16]
  reg [255:0] mem_592; // @[Ram.scala 16:16]
  reg [255:0] mem_593; // @[Ram.scala 16:16]
  reg [255:0] mem_594; // @[Ram.scala 16:16]
  reg [255:0] mem_595; // @[Ram.scala 16:16]
  reg [255:0] mem_596; // @[Ram.scala 16:16]
  reg [255:0] mem_597; // @[Ram.scala 16:16]
  reg [255:0] mem_598; // @[Ram.scala 16:16]
  reg [255:0] mem_599; // @[Ram.scala 16:16]
  reg [255:0] mem_600; // @[Ram.scala 16:16]
  reg [255:0] mem_601; // @[Ram.scala 16:16]
  reg [255:0] mem_602; // @[Ram.scala 16:16]
  reg [255:0] mem_603; // @[Ram.scala 16:16]
  reg [255:0] mem_604; // @[Ram.scala 16:16]
  reg [255:0] mem_605; // @[Ram.scala 16:16]
  reg [255:0] mem_606; // @[Ram.scala 16:16]
  reg [255:0] mem_607; // @[Ram.scala 16:16]
  reg [255:0] mem_608; // @[Ram.scala 16:16]
  reg [255:0] mem_609; // @[Ram.scala 16:16]
  reg [255:0] mem_610; // @[Ram.scala 16:16]
  reg [255:0] mem_611; // @[Ram.scala 16:16]
  reg [255:0] mem_612; // @[Ram.scala 16:16]
  reg [255:0] mem_613; // @[Ram.scala 16:16]
  reg [255:0] mem_614; // @[Ram.scala 16:16]
  reg [255:0] mem_615; // @[Ram.scala 16:16]
  reg [255:0] mem_616; // @[Ram.scala 16:16]
  reg [255:0] mem_617; // @[Ram.scala 16:16]
  reg [255:0] mem_618; // @[Ram.scala 16:16]
  reg [255:0] mem_619; // @[Ram.scala 16:16]
  reg [255:0] mem_620; // @[Ram.scala 16:16]
  reg [255:0] mem_621; // @[Ram.scala 16:16]
  reg [255:0] mem_622; // @[Ram.scala 16:16]
  reg [255:0] mem_623; // @[Ram.scala 16:16]
  reg [255:0] mem_624; // @[Ram.scala 16:16]
  reg [255:0] mem_625; // @[Ram.scala 16:16]
  reg [255:0] mem_626; // @[Ram.scala 16:16]
  reg [255:0] mem_627; // @[Ram.scala 16:16]
  reg [255:0] mem_628; // @[Ram.scala 16:16]
  reg [255:0] mem_629; // @[Ram.scala 16:16]
  reg [255:0] mem_630; // @[Ram.scala 16:16]
  reg [255:0] mem_631; // @[Ram.scala 16:16]
  reg [255:0] mem_632; // @[Ram.scala 16:16]
  reg [255:0] mem_633; // @[Ram.scala 16:16]
  reg [255:0] mem_634; // @[Ram.scala 16:16]
  reg [255:0] mem_635; // @[Ram.scala 16:16]
  reg [255:0] mem_636; // @[Ram.scala 16:16]
  reg [255:0] mem_637; // @[Ram.scala 16:16]
  reg [255:0] mem_638; // @[Ram.scala 16:16]
  reg [255:0] mem_639; // @[Ram.scala 16:16]
  reg [255:0] mem_640; // @[Ram.scala 16:16]
  reg [255:0] mem_641; // @[Ram.scala 16:16]
  reg [255:0] mem_642; // @[Ram.scala 16:16]
  reg [255:0] mem_643; // @[Ram.scala 16:16]
  reg [255:0] mem_644; // @[Ram.scala 16:16]
  reg [255:0] mem_645; // @[Ram.scala 16:16]
  reg [255:0] mem_646; // @[Ram.scala 16:16]
  reg [255:0] mem_647; // @[Ram.scala 16:16]
  reg [255:0] mem_648; // @[Ram.scala 16:16]
  reg [255:0] mem_649; // @[Ram.scala 16:16]
  reg [255:0] mem_650; // @[Ram.scala 16:16]
  reg [255:0] mem_651; // @[Ram.scala 16:16]
  reg [255:0] mem_652; // @[Ram.scala 16:16]
  reg [255:0] mem_653; // @[Ram.scala 16:16]
  reg [255:0] mem_654; // @[Ram.scala 16:16]
  reg [255:0] mem_655; // @[Ram.scala 16:16]
  reg [255:0] mem_656; // @[Ram.scala 16:16]
  reg [255:0] mem_657; // @[Ram.scala 16:16]
  reg [255:0] mem_658; // @[Ram.scala 16:16]
  reg [255:0] mem_659; // @[Ram.scala 16:16]
  reg [255:0] mem_660; // @[Ram.scala 16:16]
  reg [255:0] mem_661; // @[Ram.scala 16:16]
  reg [255:0] mem_662; // @[Ram.scala 16:16]
  reg [255:0] mem_663; // @[Ram.scala 16:16]
  reg [255:0] mem_664; // @[Ram.scala 16:16]
  reg [255:0] mem_665; // @[Ram.scala 16:16]
  reg [255:0] mem_666; // @[Ram.scala 16:16]
  reg [255:0] mem_667; // @[Ram.scala 16:16]
  reg [255:0] mem_668; // @[Ram.scala 16:16]
  reg [255:0] mem_669; // @[Ram.scala 16:16]
  reg [255:0] mem_670; // @[Ram.scala 16:16]
  reg [255:0] mem_671; // @[Ram.scala 16:16]
  reg [255:0] mem_672; // @[Ram.scala 16:16]
  reg [255:0] mem_673; // @[Ram.scala 16:16]
  reg [255:0] mem_674; // @[Ram.scala 16:16]
  reg [255:0] mem_675; // @[Ram.scala 16:16]
  reg [255:0] mem_676; // @[Ram.scala 16:16]
  reg [255:0] mem_677; // @[Ram.scala 16:16]
  reg [255:0] mem_678; // @[Ram.scala 16:16]
  reg [255:0] mem_679; // @[Ram.scala 16:16]
  reg [255:0] mem_680; // @[Ram.scala 16:16]
  reg [255:0] mem_681; // @[Ram.scala 16:16]
  reg [255:0] mem_682; // @[Ram.scala 16:16]
  reg [255:0] mem_683; // @[Ram.scala 16:16]
  reg [255:0] mem_684; // @[Ram.scala 16:16]
  reg [255:0] mem_685; // @[Ram.scala 16:16]
  reg [255:0] mem_686; // @[Ram.scala 16:16]
  reg [255:0] mem_687; // @[Ram.scala 16:16]
  reg [255:0] mem_688; // @[Ram.scala 16:16]
  reg [255:0] mem_689; // @[Ram.scala 16:16]
  reg [255:0] mem_690; // @[Ram.scala 16:16]
  reg [255:0] mem_691; // @[Ram.scala 16:16]
  reg [255:0] mem_692; // @[Ram.scala 16:16]
  reg [255:0] mem_693; // @[Ram.scala 16:16]
  reg [255:0] mem_694; // @[Ram.scala 16:16]
  reg [255:0] mem_695; // @[Ram.scala 16:16]
  reg [255:0] mem_696; // @[Ram.scala 16:16]
  reg [255:0] mem_697; // @[Ram.scala 16:16]
  reg [255:0] mem_698; // @[Ram.scala 16:16]
  reg [255:0] mem_699; // @[Ram.scala 16:16]
  reg [255:0] mem_700; // @[Ram.scala 16:16]
  reg [255:0] mem_701; // @[Ram.scala 16:16]
  reg [255:0] mem_702; // @[Ram.scala 16:16]
  reg [255:0] mem_703; // @[Ram.scala 16:16]
  reg [255:0] mem_704; // @[Ram.scala 16:16]
  reg [255:0] mem_705; // @[Ram.scala 16:16]
  reg [255:0] mem_706; // @[Ram.scala 16:16]
  reg [255:0] mem_707; // @[Ram.scala 16:16]
  reg [255:0] mem_708; // @[Ram.scala 16:16]
  reg [255:0] mem_709; // @[Ram.scala 16:16]
  reg [255:0] mem_710; // @[Ram.scala 16:16]
  reg [255:0] mem_711; // @[Ram.scala 16:16]
  reg [255:0] mem_712; // @[Ram.scala 16:16]
  reg [255:0] mem_713; // @[Ram.scala 16:16]
  reg [255:0] mem_714; // @[Ram.scala 16:16]
  reg [255:0] mem_715; // @[Ram.scala 16:16]
  reg [255:0] mem_716; // @[Ram.scala 16:16]
  reg [255:0] mem_717; // @[Ram.scala 16:16]
  reg [255:0] mem_718; // @[Ram.scala 16:16]
  reg [255:0] mem_719; // @[Ram.scala 16:16]
  reg [255:0] mem_720; // @[Ram.scala 16:16]
  reg [255:0] mem_721; // @[Ram.scala 16:16]
  reg [255:0] mem_722; // @[Ram.scala 16:16]
  reg [255:0] mem_723; // @[Ram.scala 16:16]
  reg [255:0] mem_724; // @[Ram.scala 16:16]
  reg [255:0] mem_725; // @[Ram.scala 16:16]
  reg [255:0] mem_726; // @[Ram.scala 16:16]
  reg [255:0] mem_727; // @[Ram.scala 16:16]
  reg [255:0] mem_728; // @[Ram.scala 16:16]
  reg [255:0] mem_729; // @[Ram.scala 16:16]
  reg [255:0] mem_730; // @[Ram.scala 16:16]
  reg [255:0] mem_731; // @[Ram.scala 16:16]
  reg [255:0] mem_732; // @[Ram.scala 16:16]
  reg [255:0] mem_733; // @[Ram.scala 16:16]
  reg [255:0] mem_734; // @[Ram.scala 16:16]
  reg [255:0] mem_735; // @[Ram.scala 16:16]
  reg [255:0] mem_736; // @[Ram.scala 16:16]
  reg [255:0] mem_737; // @[Ram.scala 16:16]
  reg [255:0] mem_738; // @[Ram.scala 16:16]
  reg [255:0] mem_739; // @[Ram.scala 16:16]
  reg [255:0] mem_740; // @[Ram.scala 16:16]
  reg [255:0] mem_741; // @[Ram.scala 16:16]
  reg [255:0] mem_742; // @[Ram.scala 16:16]
  reg [255:0] mem_743; // @[Ram.scala 16:16]
  reg [255:0] mem_744; // @[Ram.scala 16:16]
  reg [255:0] mem_745; // @[Ram.scala 16:16]
  reg [255:0] mem_746; // @[Ram.scala 16:16]
  reg [255:0] mem_747; // @[Ram.scala 16:16]
  reg [255:0] mem_748; // @[Ram.scala 16:16]
  reg [255:0] mem_749; // @[Ram.scala 16:16]
  reg [255:0] mem_750; // @[Ram.scala 16:16]
  reg [255:0] mem_751; // @[Ram.scala 16:16]
  reg [255:0] mem_752; // @[Ram.scala 16:16]
  reg [255:0] mem_753; // @[Ram.scala 16:16]
  reg [255:0] mem_754; // @[Ram.scala 16:16]
  reg [255:0] mem_755; // @[Ram.scala 16:16]
  reg [255:0] mem_756; // @[Ram.scala 16:16]
  reg [255:0] mem_757; // @[Ram.scala 16:16]
  reg [255:0] mem_758; // @[Ram.scala 16:16]
  reg [255:0] mem_759; // @[Ram.scala 16:16]
  reg [255:0] mem_760; // @[Ram.scala 16:16]
  reg [255:0] mem_761; // @[Ram.scala 16:16]
  reg [255:0] mem_762; // @[Ram.scala 16:16]
  reg [255:0] mem_763; // @[Ram.scala 16:16]
  reg [255:0] mem_764; // @[Ram.scala 16:16]
  reg [255:0] mem_765; // @[Ram.scala 16:16]
  reg [255:0] mem_766; // @[Ram.scala 16:16]
  reg [255:0] mem_767; // @[Ram.scala 16:16]
  reg [255:0] mem_768; // @[Ram.scala 16:16]
  reg [255:0] mem_769; // @[Ram.scala 16:16]
  reg [255:0] mem_770; // @[Ram.scala 16:16]
  reg [255:0] mem_771; // @[Ram.scala 16:16]
  reg [255:0] mem_772; // @[Ram.scala 16:16]
  reg [255:0] mem_773; // @[Ram.scala 16:16]
  reg [255:0] mem_774; // @[Ram.scala 16:16]
  reg [255:0] mem_775; // @[Ram.scala 16:16]
  reg [255:0] mem_776; // @[Ram.scala 16:16]
  reg [255:0] mem_777; // @[Ram.scala 16:16]
  reg [255:0] mem_778; // @[Ram.scala 16:16]
  reg [255:0] mem_779; // @[Ram.scala 16:16]
  reg [255:0] mem_780; // @[Ram.scala 16:16]
  reg [255:0] mem_781; // @[Ram.scala 16:16]
  reg [255:0] mem_782; // @[Ram.scala 16:16]
  reg [255:0] mem_783; // @[Ram.scala 16:16]
  reg [255:0] mem_784; // @[Ram.scala 16:16]
  reg [255:0] mem_785; // @[Ram.scala 16:16]
  reg [255:0] mem_786; // @[Ram.scala 16:16]
  reg [255:0] mem_787; // @[Ram.scala 16:16]
  reg [255:0] mem_788; // @[Ram.scala 16:16]
  reg [255:0] mem_789; // @[Ram.scala 16:16]
  reg [255:0] mem_790; // @[Ram.scala 16:16]
  reg [255:0] mem_791; // @[Ram.scala 16:16]
  reg [255:0] mem_792; // @[Ram.scala 16:16]
  reg [255:0] mem_793; // @[Ram.scala 16:16]
  reg [255:0] mem_794; // @[Ram.scala 16:16]
  reg [255:0] mem_795; // @[Ram.scala 16:16]
  reg [255:0] mem_796; // @[Ram.scala 16:16]
  reg [255:0] mem_797; // @[Ram.scala 16:16]
  reg [255:0] mem_798; // @[Ram.scala 16:16]
  reg [255:0] mem_799; // @[Ram.scala 16:16]
  reg [255:0] mem_800; // @[Ram.scala 16:16]
  reg [255:0] mem_801; // @[Ram.scala 16:16]
  reg [255:0] mem_802; // @[Ram.scala 16:16]
  reg [255:0] mem_803; // @[Ram.scala 16:16]
  reg [255:0] mem_804; // @[Ram.scala 16:16]
  reg [255:0] mem_805; // @[Ram.scala 16:16]
  reg [255:0] mem_806; // @[Ram.scala 16:16]
  reg [255:0] mem_807; // @[Ram.scala 16:16]
  reg [255:0] mem_808; // @[Ram.scala 16:16]
  reg [255:0] mem_809; // @[Ram.scala 16:16]
  reg [255:0] mem_810; // @[Ram.scala 16:16]
  reg [255:0] mem_811; // @[Ram.scala 16:16]
  reg [255:0] mem_812; // @[Ram.scala 16:16]
  reg [255:0] mem_813; // @[Ram.scala 16:16]
  reg [255:0] mem_814; // @[Ram.scala 16:16]
  reg [255:0] mem_815; // @[Ram.scala 16:16]
  reg [255:0] mem_816; // @[Ram.scala 16:16]
  reg [255:0] mem_817; // @[Ram.scala 16:16]
  reg [255:0] mem_818; // @[Ram.scala 16:16]
  reg [255:0] mem_819; // @[Ram.scala 16:16]
  reg [255:0] mem_820; // @[Ram.scala 16:16]
  reg [255:0] mem_821; // @[Ram.scala 16:16]
  reg [255:0] mem_822; // @[Ram.scala 16:16]
  reg [255:0] mem_823; // @[Ram.scala 16:16]
  reg [255:0] mem_824; // @[Ram.scala 16:16]
  reg [255:0] mem_825; // @[Ram.scala 16:16]
  reg [255:0] mem_826; // @[Ram.scala 16:16]
  reg [255:0] mem_827; // @[Ram.scala 16:16]
  reg [255:0] mem_828; // @[Ram.scala 16:16]
  reg [255:0] mem_829; // @[Ram.scala 16:16]
  reg [255:0] mem_830; // @[Ram.scala 16:16]
  reg [255:0] mem_831; // @[Ram.scala 16:16]
  reg [255:0] mem_832; // @[Ram.scala 16:16]
  reg [255:0] mem_833; // @[Ram.scala 16:16]
  reg [255:0] mem_834; // @[Ram.scala 16:16]
  reg [255:0] mem_835; // @[Ram.scala 16:16]
  reg [255:0] mem_836; // @[Ram.scala 16:16]
  reg [255:0] mem_837; // @[Ram.scala 16:16]
  reg [255:0] mem_838; // @[Ram.scala 16:16]
  reg [255:0] mem_839; // @[Ram.scala 16:16]
  reg [255:0] mem_840; // @[Ram.scala 16:16]
  reg [255:0] mem_841; // @[Ram.scala 16:16]
  reg [255:0] mem_842; // @[Ram.scala 16:16]
  reg [255:0] mem_843; // @[Ram.scala 16:16]
  reg [255:0] mem_844; // @[Ram.scala 16:16]
  reg [255:0] mem_845; // @[Ram.scala 16:16]
  reg [255:0] mem_846; // @[Ram.scala 16:16]
  reg [255:0] mem_847; // @[Ram.scala 16:16]
  reg [255:0] mem_848; // @[Ram.scala 16:16]
  reg [255:0] mem_849; // @[Ram.scala 16:16]
  reg [255:0] mem_850; // @[Ram.scala 16:16]
  reg [255:0] mem_851; // @[Ram.scala 16:16]
  reg [255:0] mem_852; // @[Ram.scala 16:16]
  reg [255:0] mem_853; // @[Ram.scala 16:16]
  reg [255:0] mem_854; // @[Ram.scala 16:16]
  reg [255:0] mem_855; // @[Ram.scala 16:16]
  reg [255:0] mem_856; // @[Ram.scala 16:16]
  reg [255:0] mem_857; // @[Ram.scala 16:16]
  reg [255:0] mem_858; // @[Ram.scala 16:16]
  reg [255:0] mem_859; // @[Ram.scala 16:16]
  reg [255:0] mem_860; // @[Ram.scala 16:16]
  reg [255:0] mem_861; // @[Ram.scala 16:16]
  reg [255:0] mem_862; // @[Ram.scala 16:16]
  reg [255:0] mem_863; // @[Ram.scala 16:16]
  reg [255:0] mem_864; // @[Ram.scala 16:16]
  reg [255:0] mem_865; // @[Ram.scala 16:16]
  reg [255:0] mem_866; // @[Ram.scala 16:16]
  reg [255:0] mem_867; // @[Ram.scala 16:16]
  reg [255:0] mem_868; // @[Ram.scala 16:16]
  reg [255:0] mem_869; // @[Ram.scala 16:16]
  reg [255:0] mem_870; // @[Ram.scala 16:16]
  reg [255:0] mem_871; // @[Ram.scala 16:16]
  reg [255:0] mem_872; // @[Ram.scala 16:16]
  reg [255:0] mem_873; // @[Ram.scala 16:16]
  reg [255:0] mem_874; // @[Ram.scala 16:16]
  reg [255:0] mem_875; // @[Ram.scala 16:16]
  reg [255:0] mem_876; // @[Ram.scala 16:16]
  reg [255:0] mem_877; // @[Ram.scala 16:16]
  reg [255:0] mem_878; // @[Ram.scala 16:16]
  reg [255:0] mem_879; // @[Ram.scala 16:16]
  reg [255:0] mem_880; // @[Ram.scala 16:16]
  reg [255:0] mem_881; // @[Ram.scala 16:16]
  reg [255:0] mem_882; // @[Ram.scala 16:16]
  reg [255:0] mem_883; // @[Ram.scala 16:16]
  reg [255:0] mem_884; // @[Ram.scala 16:16]
  reg [255:0] mem_885; // @[Ram.scala 16:16]
  reg [255:0] mem_886; // @[Ram.scala 16:16]
  reg [255:0] mem_887; // @[Ram.scala 16:16]
  reg [255:0] mem_888; // @[Ram.scala 16:16]
  reg [255:0] mem_889; // @[Ram.scala 16:16]
  reg [255:0] mem_890; // @[Ram.scala 16:16]
  reg [255:0] mem_891; // @[Ram.scala 16:16]
  reg [255:0] mem_892; // @[Ram.scala 16:16]
  reg [255:0] mem_893; // @[Ram.scala 16:16]
  reg [255:0] mem_894; // @[Ram.scala 16:16]
  reg [255:0] mem_895; // @[Ram.scala 16:16]
  reg [255:0] mem_896; // @[Ram.scala 16:16]
  reg [255:0] mem_897; // @[Ram.scala 16:16]
  reg [255:0] mem_898; // @[Ram.scala 16:16]
  reg [255:0] mem_899; // @[Ram.scala 16:16]
  reg [255:0] mem_900; // @[Ram.scala 16:16]
  reg [255:0] mem_901; // @[Ram.scala 16:16]
  reg [255:0] mem_902; // @[Ram.scala 16:16]
  reg [255:0] mem_903; // @[Ram.scala 16:16]
  reg [255:0] mem_904; // @[Ram.scala 16:16]
  reg [255:0] mem_905; // @[Ram.scala 16:16]
  reg [255:0] mem_906; // @[Ram.scala 16:16]
  reg [255:0] mem_907; // @[Ram.scala 16:16]
  reg [255:0] mem_908; // @[Ram.scala 16:16]
  reg [255:0] mem_909; // @[Ram.scala 16:16]
  reg [255:0] mem_910; // @[Ram.scala 16:16]
  reg [255:0] mem_911; // @[Ram.scala 16:16]
  reg [255:0] mem_912; // @[Ram.scala 16:16]
  reg [255:0] mem_913; // @[Ram.scala 16:16]
  reg [255:0] mem_914; // @[Ram.scala 16:16]
  reg [255:0] mem_915; // @[Ram.scala 16:16]
  reg [255:0] mem_916; // @[Ram.scala 16:16]
  reg [255:0] mem_917; // @[Ram.scala 16:16]
  reg [255:0] mem_918; // @[Ram.scala 16:16]
  reg [255:0] mem_919; // @[Ram.scala 16:16]
  reg [255:0] mem_920; // @[Ram.scala 16:16]
  reg [255:0] mem_921; // @[Ram.scala 16:16]
  reg [255:0] mem_922; // @[Ram.scala 16:16]
  reg [255:0] mem_923; // @[Ram.scala 16:16]
  reg [255:0] mem_924; // @[Ram.scala 16:16]
  reg [255:0] mem_925; // @[Ram.scala 16:16]
  reg [255:0] mem_926; // @[Ram.scala 16:16]
  reg [255:0] mem_927; // @[Ram.scala 16:16]
  reg [255:0] mem_928; // @[Ram.scala 16:16]
  reg [255:0] mem_929; // @[Ram.scala 16:16]
  reg [255:0] mem_930; // @[Ram.scala 16:16]
  reg [255:0] mem_931; // @[Ram.scala 16:16]
  reg [255:0] mem_932; // @[Ram.scala 16:16]
  reg [255:0] mem_933; // @[Ram.scala 16:16]
  reg [255:0] mem_934; // @[Ram.scala 16:16]
  reg [255:0] mem_935; // @[Ram.scala 16:16]
  reg [255:0] mem_936; // @[Ram.scala 16:16]
  reg [255:0] mem_937; // @[Ram.scala 16:16]
  reg [255:0] mem_938; // @[Ram.scala 16:16]
  reg [255:0] mem_939; // @[Ram.scala 16:16]
  reg [255:0] mem_940; // @[Ram.scala 16:16]
  reg [255:0] mem_941; // @[Ram.scala 16:16]
  reg [255:0] mem_942; // @[Ram.scala 16:16]
  reg [255:0] mem_943; // @[Ram.scala 16:16]
  reg [255:0] mem_944; // @[Ram.scala 16:16]
  reg [255:0] mem_945; // @[Ram.scala 16:16]
  reg [255:0] mem_946; // @[Ram.scala 16:16]
  reg [255:0] mem_947; // @[Ram.scala 16:16]
  reg [255:0] mem_948; // @[Ram.scala 16:16]
  reg [255:0] mem_949; // @[Ram.scala 16:16]
  reg [255:0] mem_950; // @[Ram.scala 16:16]
  reg [255:0] mem_951; // @[Ram.scala 16:16]
  reg [255:0] mem_952; // @[Ram.scala 16:16]
  reg [255:0] mem_953; // @[Ram.scala 16:16]
  reg [255:0] mem_954; // @[Ram.scala 16:16]
  reg [255:0] mem_955; // @[Ram.scala 16:16]
  reg [255:0] mem_956; // @[Ram.scala 16:16]
  reg [255:0] mem_957; // @[Ram.scala 16:16]
  reg [255:0] mem_958; // @[Ram.scala 16:16]
  reg [255:0] mem_959; // @[Ram.scala 16:16]
  reg [255:0] mem_960; // @[Ram.scala 16:16]
  reg [255:0] mem_961; // @[Ram.scala 16:16]
  reg [255:0] mem_962; // @[Ram.scala 16:16]
  reg [255:0] mem_963; // @[Ram.scala 16:16]
  reg [255:0] mem_964; // @[Ram.scala 16:16]
  reg [255:0] mem_965; // @[Ram.scala 16:16]
  reg [255:0] mem_966; // @[Ram.scala 16:16]
  reg [255:0] mem_967; // @[Ram.scala 16:16]
  reg [255:0] mem_968; // @[Ram.scala 16:16]
  reg [255:0] mem_969; // @[Ram.scala 16:16]
  reg [255:0] mem_970; // @[Ram.scala 16:16]
  reg [255:0] mem_971; // @[Ram.scala 16:16]
  reg [255:0] mem_972; // @[Ram.scala 16:16]
  reg [255:0] mem_973; // @[Ram.scala 16:16]
  reg [255:0] mem_974; // @[Ram.scala 16:16]
  reg [255:0] mem_975; // @[Ram.scala 16:16]
  reg [255:0] mem_976; // @[Ram.scala 16:16]
  reg [255:0] mem_977; // @[Ram.scala 16:16]
  reg [255:0] mem_978; // @[Ram.scala 16:16]
  reg [255:0] mem_979; // @[Ram.scala 16:16]
  reg [255:0] mem_980; // @[Ram.scala 16:16]
  reg [255:0] mem_981; // @[Ram.scala 16:16]
  reg [255:0] mem_982; // @[Ram.scala 16:16]
  reg [255:0] mem_983; // @[Ram.scala 16:16]
  reg [255:0] mem_984; // @[Ram.scala 16:16]
  reg [255:0] mem_985; // @[Ram.scala 16:16]
  reg [255:0] mem_986; // @[Ram.scala 16:16]
  reg [255:0] mem_987; // @[Ram.scala 16:16]
  reg [255:0] mem_988; // @[Ram.scala 16:16]
  reg [255:0] mem_989; // @[Ram.scala 16:16]
  reg [255:0] mem_990; // @[Ram.scala 16:16]
  reg [255:0] mem_991; // @[Ram.scala 16:16]
  reg [255:0] mem_992; // @[Ram.scala 16:16]
  reg [255:0] mem_993; // @[Ram.scala 16:16]
  reg [255:0] mem_994; // @[Ram.scala 16:16]
  reg [255:0] mem_995; // @[Ram.scala 16:16]
  reg [255:0] mem_996; // @[Ram.scala 16:16]
  reg [255:0] mem_997; // @[Ram.scala 16:16]
  reg [255:0] mem_998; // @[Ram.scala 16:16]
  reg [255:0] mem_999; // @[Ram.scala 16:16]
  reg [255:0] mem_1000; // @[Ram.scala 16:16]
  reg [255:0] mem_1001; // @[Ram.scala 16:16]
  reg [255:0] mem_1002; // @[Ram.scala 16:16]
  reg [255:0] mem_1003; // @[Ram.scala 16:16]
  reg [255:0] mem_1004; // @[Ram.scala 16:16]
  reg [255:0] mem_1005; // @[Ram.scala 16:16]
  reg [255:0] mem_1006; // @[Ram.scala 16:16]
  reg [255:0] mem_1007; // @[Ram.scala 16:16]
  reg [255:0] mem_1008; // @[Ram.scala 16:16]
  reg [255:0] mem_1009; // @[Ram.scala 16:16]
  reg [255:0] mem_1010; // @[Ram.scala 16:16]
  reg [255:0] mem_1011; // @[Ram.scala 16:16]
  reg [255:0] mem_1012; // @[Ram.scala 16:16]
  reg [255:0] mem_1013; // @[Ram.scala 16:16]
  reg [255:0] mem_1014; // @[Ram.scala 16:16]
  reg [255:0] mem_1015; // @[Ram.scala 16:16]
  reg [255:0] mem_1016; // @[Ram.scala 16:16]
  reg [255:0] mem_1017; // @[Ram.scala 16:16]
  reg [255:0] mem_1018; // @[Ram.scala 16:16]
  reg [255:0] mem_1019; // @[Ram.scala 16:16]
  reg [255:0] mem_1020; // @[Ram.scala 16:16]
  reg [255:0] mem_1021; // @[Ram.scala 16:16]
  reg [255:0] mem_1022; // @[Ram.scala 16:16]
  reg [255:0] mem_1023; // @[Ram.scala 16:16]
  wire [255:0] _GEN_1025 = 10'h1 == io_addr ? mem_1 : mem_0; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1026 = 10'h2 == io_addr ? mem_2 : _GEN_1025; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1027 = 10'h3 == io_addr ? mem_3 : _GEN_1026; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1028 = 10'h4 == io_addr ? mem_4 : _GEN_1027; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1029 = 10'h5 == io_addr ? mem_5 : _GEN_1028; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1030 = 10'h6 == io_addr ? mem_6 : _GEN_1029; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1031 = 10'h7 == io_addr ? mem_7 : _GEN_1030; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1032 = 10'h8 == io_addr ? mem_8 : _GEN_1031; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1033 = 10'h9 == io_addr ? mem_9 : _GEN_1032; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1034 = 10'ha == io_addr ? mem_10 : _GEN_1033; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1035 = 10'hb == io_addr ? mem_11 : _GEN_1034; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1036 = 10'hc == io_addr ? mem_12 : _GEN_1035; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1037 = 10'hd == io_addr ? mem_13 : _GEN_1036; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1038 = 10'he == io_addr ? mem_14 : _GEN_1037; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1039 = 10'hf == io_addr ? mem_15 : _GEN_1038; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1040 = 10'h10 == io_addr ? mem_16 : _GEN_1039; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1041 = 10'h11 == io_addr ? mem_17 : _GEN_1040; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1042 = 10'h12 == io_addr ? mem_18 : _GEN_1041; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1043 = 10'h13 == io_addr ? mem_19 : _GEN_1042; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1044 = 10'h14 == io_addr ? mem_20 : _GEN_1043; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1045 = 10'h15 == io_addr ? mem_21 : _GEN_1044; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1046 = 10'h16 == io_addr ? mem_22 : _GEN_1045; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1047 = 10'h17 == io_addr ? mem_23 : _GEN_1046; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1048 = 10'h18 == io_addr ? mem_24 : _GEN_1047; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1049 = 10'h19 == io_addr ? mem_25 : _GEN_1048; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1050 = 10'h1a == io_addr ? mem_26 : _GEN_1049; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1051 = 10'h1b == io_addr ? mem_27 : _GEN_1050; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1052 = 10'h1c == io_addr ? mem_28 : _GEN_1051; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1053 = 10'h1d == io_addr ? mem_29 : _GEN_1052; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1054 = 10'h1e == io_addr ? mem_30 : _GEN_1053; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1055 = 10'h1f == io_addr ? mem_31 : _GEN_1054; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1056 = 10'h20 == io_addr ? mem_32 : _GEN_1055; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1057 = 10'h21 == io_addr ? mem_33 : _GEN_1056; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1058 = 10'h22 == io_addr ? mem_34 : _GEN_1057; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1059 = 10'h23 == io_addr ? mem_35 : _GEN_1058; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1060 = 10'h24 == io_addr ? mem_36 : _GEN_1059; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1061 = 10'h25 == io_addr ? mem_37 : _GEN_1060; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1062 = 10'h26 == io_addr ? mem_38 : _GEN_1061; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1063 = 10'h27 == io_addr ? mem_39 : _GEN_1062; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1064 = 10'h28 == io_addr ? mem_40 : _GEN_1063; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1065 = 10'h29 == io_addr ? mem_41 : _GEN_1064; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1066 = 10'h2a == io_addr ? mem_42 : _GEN_1065; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1067 = 10'h2b == io_addr ? mem_43 : _GEN_1066; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1068 = 10'h2c == io_addr ? mem_44 : _GEN_1067; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1069 = 10'h2d == io_addr ? mem_45 : _GEN_1068; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1070 = 10'h2e == io_addr ? mem_46 : _GEN_1069; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1071 = 10'h2f == io_addr ? mem_47 : _GEN_1070; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1072 = 10'h30 == io_addr ? mem_48 : _GEN_1071; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1073 = 10'h31 == io_addr ? mem_49 : _GEN_1072; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1074 = 10'h32 == io_addr ? mem_50 : _GEN_1073; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1075 = 10'h33 == io_addr ? mem_51 : _GEN_1074; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1076 = 10'h34 == io_addr ? mem_52 : _GEN_1075; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1077 = 10'h35 == io_addr ? mem_53 : _GEN_1076; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1078 = 10'h36 == io_addr ? mem_54 : _GEN_1077; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1079 = 10'h37 == io_addr ? mem_55 : _GEN_1078; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1080 = 10'h38 == io_addr ? mem_56 : _GEN_1079; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1081 = 10'h39 == io_addr ? mem_57 : _GEN_1080; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1082 = 10'h3a == io_addr ? mem_58 : _GEN_1081; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1083 = 10'h3b == io_addr ? mem_59 : _GEN_1082; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1084 = 10'h3c == io_addr ? mem_60 : _GEN_1083; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1085 = 10'h3d == io_addr ? mem_61 : _GEN_1084; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1086 = 10'h3e == io_addr ? mem_62 : _GEN_1085; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1087 = 10'h3f == io_addr ? mem_63 : _GEN_1086; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1088 = 10'h40 == io_addr ? mem_64 : _GEN_1087; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1089 = 10'h41 == io_addr ? mem_65 : _GEN_1088; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1090 = 10'h42 == io_addr ? mem_66 : _GEN_1089; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1091 = 10'h43 == io_addr ? mem_67 : _GEN_1090; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1092 = 10'h44 == io_addr ? mem_68 : _GEN_1091; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1093 = 10'h45 == io_addr ? mem_69 : _GEN_1092; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1094 = 10'h46 == io_addr ? mem_70 : _GEN_1093; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1095 = 10'h47 == io_addr ? mem_71 : _GEN_1094; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1096 = 10'h48 == io_addr ? mem_72 : _GEN_1095; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1097 = 10'h49 == io_addr ? mem_73 : _GEN_1096; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1098 = 10'h4a == io_addr ? mem_74 : _GEN_1097; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1099 = 10'h4b == io_addr ? mem_75 : _GEN_1098; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1100 = 10'h4c == io_addr ? mem_76 : _GEN_1099; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1101 = 10'h4d == io_addr ? mem_77 : _GEN_1100; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1102 = 10'h4e == io_addr ? mem_78 : _GEN_1101; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1103 = 10'h4f == io_addr ? mem_79 : _GEN_1102; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1104 = 10'h50 == io_addr ? mem_80 : _GEN_1103; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1105 = 10'h51 == io_addr ? mem_81 : _GEN_1104; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1106 = 10'h52 == io_addr ? mem_82 : _GEN_1105; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1107 = 10'h53 == io_addr ? mem_83 : _GEN_1106; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1108 = 10'h54 == io_addr ? mem_84 : _GEN_1107; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1109 = 10'h55 == io_addr ? mem_85 : _GEN_1108; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1110 = 10'h56 == io_addr ? mem_86 : _GEN_1109; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1111 = 10'h57 == io_addr ? mem_87 : _GEN_1110; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1112 = 10'h58 == io_addr ? mem_88 : _GEN_1111; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1113 = 10'h59 == io_addr ? mem_89 : _GEN_1112; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1114 = 10'h5a == io_addr ? mem_90 : _GEN_1113; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1115 = 10'h5b == io_addr ? mem_91 : _GEN_1114; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1116 = 10'h5c == io_addr ? mem_92 : _GEN_1115; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1117 = 10'h5d == io_addr ? mem_93 : _GEN_1116; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1118 = 10'h5e == io_addr ? mem_94 : _GEN_1117; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1119 = 10'h5f == io_addr ? mem_95 : _GEN_1118; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1120 = 10'h60 == io_addr ? mem_96 : _GEN_1119; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1121 = 10'h61 == io_addr ? mem_97 : _GEN_1120; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1122 = 10'h62 == io_addr ? mem_98 : _GEN_1121; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1123 = 10'h63 == io_addr ? mem_99 : _GEN_1122; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1124 = 10'h64 == io_addr ? mem_100 : _GEN_1123; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1125 = 10'h65 == io_addr ? mem_101 : _GEN_1124; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1126 = 10'h66 == io_addr ? mem_102 : _GEN_1125; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1127 = 10'h67 == io_addr ? mem_103 : _GEN_1126; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1128 = 10'h68 == io_addr ? mem_104 : _GEN_1127; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1129 = 10'h69 == io_addr ? mem_105 : _GEN_1128; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1130 = 10'h6a == io_addr ? mem_106 : _GEN_1129; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1131 = 10'h6b == io_addr ? mem_107 : _GEN_1130; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1132 = 10'h6c == io_addr ? mem_108 : _GEN_1131; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1133 = 10'h6d == io_addr ? mem_109 : _GEN_1132; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1134 = 10'h6e == io_addr ? mem_110 : _GEN_1133; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1135 = 10'h6f == io_addr ? mem_111 : _GEN_1134; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1136 = 10'h70 == io_addr ? mem_112 : _GEN_1135; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1137 = 10'h71 == io_addr ? mem_113 : _GEN_1136; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1138 = 10'h72 == io_addr ? mem_114 : _GEN_1137; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1139 = 10'h73 == io_addr ? mem_115 : _GEN_1138; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1140 = 10'h74 == io_addr ? mem_116 : _GEN_1139; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1141 = 10'h75 == io_addr ? mem_117 : _GEN_1140; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1142 = 10'h76 == io_addr ? mem_118 : _GEN_1141; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1143 = 10'h77 == io_addr ? mem_119 : _GEN_1142; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1144 = 10'h78 == io_addr ? mem_120 : _GEN_1143; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1145 = 10'h79 == io_addr ? mem_121 : _GEN_1144; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1146 = 10'h7a == io_addr ? mem_122 : _GEN_1145; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1147 = 10'h7b == io_addr ? mem_123 : _GEN_1146; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1148 = 10'h7c == io_addr ? mem_124 : _GEN_1147; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1149 = 10'h7d == io_addr ? mem_125 : _GEN_1148; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1150 = 10'h7e == io_addr ? mem_126 : _GEN_1149; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1151 = 10'h7f == io_addr ? mem_127 : _GEN_1150; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1152 = 10'h80 == io_addr ? mem_128 : _GEN_1151; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1153 = 10'h81 == io_addr ? mem_129 : _GEN_1152; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1154 = 10'h82 == io_addr ? mem_130 : _GEN_1153; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1155 = 10'h83 == io_addr ? mem_131 : _GEN_1154; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1156 = 10'h84 == io_addr ? mem_132 : _GEN_1155; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1157 = 10'h85 == io_addr ? mem_133 : _GEN_1156; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1158 = 10'h86 == io_addr ? mem_134 : _GEN_1157; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1159 = 10'h87 == io_addr ? mem_135 : _GEN_1158; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1160 = 10'h88 == io_addr ? mem_136 : _GEN_1159; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1161 = 10'h89 == io_addr ? mem_137 : _GEN_1160; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1162 = 10'h8a == io_addr ? mem_138 : _GEN_1161; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1163 = 10'h8b == io_addr ? mem_139 : _GEN_1162; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1164 = 10'h8c == io_addr ? mem_140 : _GEN_1163; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1165 = 10'h8d == io_addr ? mem_141 : _GEN_1164; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1166 = 10'h8e == io_addr ? mem_142 : _GEN_1165; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1167 = 10'h8f == io_addr ? mem_143 : _GEN_1166; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1168 = 10'h90 == io_addr ? mem_144 : _GEN_1167; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1169 = 10'h91 == io_addr ? mem_145 : _GEN_1168; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1170 = 10'h92 == io_addr ? mem_146 : _GEN_1169; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1171 = 10'h93 == io_addr ? mem_147 : _GEN_1170; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1172 = 10'h94 == io_addr ? mem_148 : _GEN_1171; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1173 = 10'h95 == io_addr ? mem_149 : _GEN_1172; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1174 = 10'h96 == io_addr ? mem_150 : _GEN_1173; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1175 = 10'h97 == io_addr ? mem_151 : _GEN_1174; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1176 = 10'h98 == io_addr ? mem_152 : _GEN_1175; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1177 = 10'h99 == io_addr ? mem_153 : _GEN_1176; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1178 = 10'h9a == io_addr ? mem_154 : _GEN_1177; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1179 = 10'h9b == io_addr ? mem_155 : _GEN_1178; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1180 = 10'h9c == io_addr ? mem_156 : _GEN_1179; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1181 = 10'h9d == io_addr ? mem_157 : _GEN_1180; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1182 = 10'h9e == io_addr ? mem_158 : _GEN_1181; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1183 = 10'h9f == io_addr ? mem_159 : _GEN_1182; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1184 = 10'ha0 == io_addr ? mem_160 : _GEN_1183; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1185 = 10'ha1 == io_addr ? mem_161 : _GEN_1184; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1186 = 10'ha2 == io_addr ? mem_162 : _GEN_1185; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1187 = 10'ha3 == io_addr ? mem_163 : _GEN_1186; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1188 = 10'ha4 == io_addr ? mem_164 : _GEN_1187; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1189 = 10'ha5 == io_addr ? mem_165 : _GEN_1188; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1190 = 10'ha6 == io_addr ? mem_166 : _GEN_1189; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1191 = 10'ha7 == io_addr ? mem_167 : _GEN_1190; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1192 = 10'ha8 == io_addr ? mem_168 : _GEN_1191; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1193 = 10'ha9 == io_addr ? mem_169 : _GEN_1192; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1194 = 10'haa == io_addr ? mem_170 : _GEN_1193; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1195 = 10'hab == io_addr ? mem_171 : _GEN_1194; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1196 = 10'hac == io_addr ? mem_172 : _GEN_1195; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1197 = 10'had == io_addr ? mem_173 : _GEN_1196; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1198 = 10'hae == io_addr ? mem_174 : _GEN_1197; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1199 = 10'haf == io_addr ? mem_175 : _GEN_1198; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1200 = 10'hb0 == io_addr ? mem_176 : _GEN_1199; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1201 = 10'hb1 == io_addr ? mem_177 : _GEN_1200; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1202 = 10'hb2 == io_addr ? mem_178 : _GEN_1201; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1203 = 10'hb3 == io_addr ? mem_179 : _GEN_1202; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1204 = 10'hb4 == io_addr ? mem_180 : _GEN_1203; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1205 = 10'hb5 == io_addr ? mem_181 : _GEN_1204; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1206 = 10'hb6 == io_addr ? mem_182 : _GEN_1205; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1207 = 10'hb7 == io_addr ? mem_183 : _GEN_1206; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1208 = 10'hb8 == io_addr ? mem_184 : _GEN_1207; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1209 = 10'hb9 == io_addr ? mem_185 : _GEN_1208; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1210 = 10'hba == io_addr ? mem_186 : _GEN_1209; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1211 = 10'hbb == io_addr ? mem_187 : _GEN_1210; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1212 = 10'hbc == io_addr ? mem_188 : _GEN_1211; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1213 = 10'hbd == io_addr ? mem_189 : _GEN_1212; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1214 = 10'hbe == io_addr ? mem_190 : _GEN_1213; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1215 = 10'hbf == io_addr ? mem_191 : _GEN_1214; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1216 = 10'hc0 == io_addr ? mem_192 : _GEN_1215; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1217 = 10'hc1 == io_addr ? mem_193 : _GEN_1216; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1218 = 10'hc2 == io_addr ? mem_194 : _GEN_1217; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1219 = 10'hc3 == io_addr ? mem_195 : _GEN_1218; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1220 = 10'hc4 == io_addr ? mem_196 : _GEN_1219; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1221 = 10'hc5 == io_addr ? mem_197 : _GEN_1220; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1222 = 10'hc6 == io_addr ? mem_198 : _GEN_1221; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1223 = 10'hc7 == io_addr ? mem_199 : _GEN_1222; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1224 = 10'hc8 == io_addr ? mem_200 : _GEN_1223; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1225 = 10'hc9 == io_addr ? mem_201 : _GEN_1224; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1226 = 10'hca == io_addr ? mem_202 : _GEN_1225; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1227 = 10'hcb == io_addr ? mem_203 : _GEN_1226; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1228 = 10'hcc == io_addr ? mem_204 : _GEN_1227; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1229 = 10'hcd == io_addr ? mem_205 : _GEN_1228; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1230 = 10'hce == io_addr ? mem_206 : _GEN_1229; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1231 = 10'hcf == io_addr ? mem_207 : _GEN_1230; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1232 = 10'hd0 == io_addr ? mem_208 : _GEN_1231; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1233 = 10'hd1 == io_addr ? mem_209 : _GEN_1232; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1234 = 10'hd2 == io_addr ? mem_210 : _GEN_1233; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1235 = 10'hd3 == io_addr ? mem_211 : _GEN_1234; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1236 = 10'hd4 == io_addr ? mem_212 : _GEN_1235; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1237 = 10'hd5 == io_addr ? mem_213 : _GEN_1236; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1238 = 10'hd6 == io_addr ? mem_214 : _GEN_1237; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1239 = 10'hd7 == io_addr ? mem_215 : _GEN_1238; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1240 = 10'hd8 == io_addr ? mem_216 : _GEN_1239; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1241 = 10'hd9 == io_addr ? mem_217 : _GEN_1240; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1242 = 10'hda == io_addr ? mem_218 : _GEN_1241; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1243 = 10'hdb == io_addr ? mem_219 : _GEN_1242; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1244 = 10'hdc == io_addr ? mem_220 : _GEN_1243; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1245 = 10'hdd == io_addr ? mem_221 : _GEN_1244; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1246 = 10'hde == io_addr ? mem_222 : _GEN_1245; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1247 = 10'hdf == io_addr ? mem_223 : _GEN_1246; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1248 = 10'he0 == io_addr ? mem_224 : _GEN_1247; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1249 = 10'he1 == io_addr ? mem_225 : _GEN_1248; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1250 = 10'he2 == io_addr ? mem_226 : _GEN_1249; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1251 = 10'he3 == io_addr ? mem_227 : _GEN_1250; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1252 = 10'he4 == io_addr ? mem_228 : _GEN_1251; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1253 = 10'he5 == io_addr ? mem_229 : _GEN_1252; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1254 = 10'he6 == io_addr ? mem_230 : _GEN_1253; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1255 = 10'he7 == io_addr ? mem_231 : _GEN_1254; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1256 = 10'he8 == io_addr ? mem_232 : _GEN_1255; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1257 = 10'he9 == io_addr ? mem_233 : _GEN_1256; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1258 = 10'hea == io_addr ? mem_234 : _GEN_1257; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1259 = 10'heb == io_addr ? mem_235 : _GEN_1258; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1260 = 10'hec == io_addr ? mem_236 : _GEN_1259; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1261 = 10'hed == io_addr ? mem_237 : _GEN_1260; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1262 = 10'hee == io_addr ? mem_238 : _GEN_1261; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1263 = 10'hef == io_addr ? mem_239 : _GEN_1262; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1264 = 10'hf0 == io_addr ? mem_240 : _GEN_1263; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1265 = 10'hf1 == io_addr ? mem_241 : _GEN_1264; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1266 = 10'hf2 == io_addr ? mem_242 : _GEN_1265; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1267 = 10'hf3 == io_addr ? mem_243 : _GEN_1266; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1268 = 10'hf4 == io_addr ? mem_244 : _GEN_1267; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1269 = 10'hf5 == io_addr ? mem_245 : _GEN_1268; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1270 = 10'hf6 == io_addr ? mem_246 : _GEN_1269; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1271 = 10'hf7 == io_addr ? mem_247 : _GEN_1270; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1272 = 10'hf8 == io_addr ? mem_248 : _GEN_1271; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1273 = 10'hf9 == io_addr ? mem_249 : _GEN_1272; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1274 = 10'hfa == io_addr ? mem_250 : _GEN_1273; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1275 = 10'hfb == io_addr ? mem_251 : _GEN_1274; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1276 = 10'hfc == io_addr ? mem_252 : _GEN_1275; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1277 = 10'hfd == io_addr ? mem_253 : _GEN_1276; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1278 = 10'hfe == io_addr ? mem_254 : _GEN_1277; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1279 = 10'hff == io_addr ? mem_255 : _GEN_1278; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1280 = 10'h100 == io_addr ? mem_256 : _GEN_1279; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1281 = 10'h101 == io_addr ? mem_257 : _GEN_1280; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1282 = 10'h102 == io_addr ? mem_258 : _GEN_1281; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1283 = 10'h103 == io_addr ? mem_259 : _GEN_1282; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1284 = 10'h104 == io_addr ? mem_260 : _GEN_1283; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1285 = 10'h105 == io_addr ? mem_261 : _GEN_1284; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1286 = 10'h106 == io_addr ? mem_262 : _GEN_1285; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1287 = 10'h107 == io_addr ? mem_263 : _GEN_1286; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1288 = 10'h108 == io_addr ? mem_264 : _GEN_1287; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1289 = 10'h109 == io_addr ? mem_265 : _GEN_1288; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1290 = 10'h10a == io_addr ? mem_266 : _GEN_1289; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1291 = 10'h10b == io_addr ? mem_267 : _GEN_1290; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1292 = 10'h10c == io_addr ? mem_268 : _GEN_1291; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1293 = 10'h10d == io_addr ? mem_269 : _GEN_1292; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1294 = 10'h10e == io_addr ? mem_270 : _GEN_1293; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1295 = 10'h10f == io_addr ? mem_271 : _GEN_1294; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1296 = 10'h110 == io_addr ? mem_272 : _GEN_1295; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1297 = 10'h111 == io_addr ? mem_273 : _GEN_1296; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1298 = 10'h112 == io_addr ? mem_274 : _GEN_1297; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1299 = 10'h113 == io_addr ? mem_275 : _GEN_1298; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1300 = 10'h114 == io_addr ? mem_276 : _GEN_1299; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1301 = 10'h115 == io_addr ? mem_277 : _GEN_1300; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1302 = 10'h116 == io_addr ? mem_278 : _GEN_1301; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1303 = 10'h117 == io_addr ? mem_279 : _GEN_1302; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1304 = 10'h118 == io_addr ? mem_280 : _GEN_1303; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1305 = 10'h119 == io_addr ? mem_281 : _GEN_1304; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1306 = 10'h11a == io_addr ? mem_282 : _GEN_1305; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1307 = 10'h11b == io_addr ? mem_283 : _GEN_1306; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1308 = 10'h11c == io_addr ? mem_284 : _GEN_1307; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1309 = 10'h11d == io_addr ? mem_285 : _GEN_1308; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1310 = 10'h11e == io_addr ? mem_286 : _GEN_1309; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1311 = 10'h11f == io_addr ? mem_287 : _GEN_1310; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1312 = 10'h120 == io_addr ? mem_288 : _GEN_1311; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1313 = 10'h121 == io_addr ? mem_289 : _GEN_1312; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1314 = 10'h122 == io_addr ? mem_290 : _GEN_1313; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1315 = 10'h123 == io_addr ? mem_291 : _GEN_1314; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1316 = 10'h124 == io_addr ? mem_292 : _GEN_1315; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1317 = 10'h125 == io_addr ? mem_293 : _GEN_1316; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1318 = 10'h126 == io_addr ? mem_294 : _GEN_1317; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1319 = 10'h127 == io_addr ? mem_295 : _GEN_1318; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1320 = 10'h128 == io_addr ? mem_296 : _GEN_1319; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1321 = 10'h129 == io_addr ? mem_297 : _GEN_1320; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1322 = 10'h12a == io_addr ? mem_298 : _GEN_1321; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1323 = 10'h12b == io_addr ? mem_299 : _GEN_1322; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1324 = 10'h12c == io_addr ? mem_300 : _GEN_1323; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1325 = 10'h12d == io_addr ? mem_301 : _GEN_1324; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1326 = 10'h12e == io_addr ? mem_302 : _GEN_1325; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1327 = 10'h12f == io_addr ? mem_303 : _GEN_1326; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1328 = 10'h130 == io_addr ? mem_304 : _GEN_1327; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1329 = 10'h131 == io_addr ? mem_305 : _GEN_1328; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1330 = 10'h132 == io_addr ? mem_306 : _GEN_1329; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1331 = 10'h133 == io_addr ? mem_307 : _GEN_1330; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1332 = 10'h134 == io_addr ? mem_308 : _GEN_1331; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1333 = 10'h135 == io_addr ? mem_309 : _GEN_1332; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1334 = 10'h136 == io_addr ? mem_310 : _GEN_1333; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1335 = 10'h137 == io_addr ? mem_311 : _GEN_1334; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1336 = 10'h138 == io_addr ? mem_312 : _GEN_1335; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1337 = 10'h139 == io_addr ? mem_313 : _GEN_1336; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1338 = 10'h13a == io_addr ? mem_314 : _GEN_1337; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1339 = 10'h13b == io_addr ? mem_315 : _GEN_1338; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1340 = 10'h13c == io_addr ? mem_316 : _GEN_1339; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1341 = 10'h13d == io_addr ? mem_317 : _GEN_1340; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1342 = 10'h13e == io_addr ? mem_318 : _GEN_1341; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1343 = 10'h13f == io_addr ? mem_319 : _GEN_1342; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1344 = 10'h140 == io_addr ? mem_320 : _GEN_1343; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1345 = 10'h141 == io_addr ? mem_321 : _GEN_1344; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1346 = 10'h142 == io_addr ? mem_322 : _GEN_1345; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1347 = 10'h143 == io_addr ? mem_323 : _GEN_1346; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1348 = 10'h144 == io_addr ? mem_324 : _GEN_1347; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1349 = 10'h145 == io_addr ? mem_325 : _GEN_1348; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1350 = 10'h146 == io_addr ? mem_326 : _GEN_1349; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1351 = 10'h147 == io_addr ? mem_327 : _GEN_1350; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1352 = 10'h148 == io_addr ? mem_328 : _GEN_1351; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1353 = 10'h149 == io_addr ? mem_329 : _GEN_1352; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1354 = 10'h14a == io_addr ? mem_330 : _GEN_1353; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1355 = 10'h14b == io_addr ? mem_331 : _GEN_1354; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1356 = 10'h14c == io_addr ? mem_332 : _GEN_1355; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1357 = 10'h14d == io_addr ? mem_333 : _GEN_1356; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1358 = 10'h14e == io_addr ? mem_334 : _GEN_1357; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1359 = 10'h14f == io_addr ? mem_335 : _GEN_1358; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1360 = 10'h150 == io_addr ? mem_336 : _GEN_1359; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1361 = 10'h151 == io_addr ? mem_337 : _GEN_1360; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1362 = 10'h152 == io_addr ? mem_338 : _GEN_1361; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1363 = 10'h153 == io_addr ? mem_339 : _GEN_1362; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1364 = 10'h154 == io_addr ? mem_340 : _GEN_1363; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1365 = 10'h155 == io_addr ? mem_341 : _GEN_1364; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1366 = 10'h156 == io_addr ? mem_342 : _GEN_1365; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1367 = 10'h157 == io_addr ? mem_343 : _GEN_1366; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1368 = 10'h158 == io_addr ? mem_344 : _GEN_1367; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1369 = 10'h159 == io_addr ? mem_345 : _GEN_1368; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1370 = 10'h15a == io_addr ? mem_346 : _GEN_1369; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1371 = 10'h15b == io_addr ? mem_347 : _GEN_1370; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1372 = 10'h15c == io_addr ? mem_348 : _GEN_1371; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1373 = 10'h15d == io_addr ? mem_349 : _GEN_1372; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1374 = 10'h15e == io_addr ? mem_350 : _GEN_1373; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1375 = 10'h15f == io_addr ? mem_351 : _GEN_1374; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1376 = 10'h160 == io_addr ? mem_352 : _GEN_1375; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1377 = 10'h161 == io_addr ? mem_353 : _GEN_1376; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1378 = 10'h162 == io_addr ? mem_354 : _GEN_1377; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1379 = 10'h163 == io_addr ? mem_355 : _GEN_1378; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1380 = 10'h164 == io_addr ? mem_356 : _GEN_1379; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1381 = 10'h165 == io_addr ? mem_357 : _GEN_1380; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1382 = 10'h166 == io_addr ? mem_358 : _GEN_1381; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1383 = 10'h167 == io_addr ? mem_359 : _GEN_1382; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1384 = 10'h168 == io_addr ? mem_360 : _GEN_1383; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1385 = 10'h169 == io_addr ? mem_361 : _GEN_1384; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1386 = 10'h16a == io_addr ? mem_362 : _GEN_1385; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1387 = 10'h16b == io_addr ? mem_363 : _GEN_1386; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1388 = 10'h16c == io_addr ? mem_364 : _GEN_1387; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1389 = 10'h16d == io_addr ? mem_365 : _GEN_1388; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1390 = 10'h16e == io_addr ? mem_366 : _GEN_1389; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1391 = 10'h16f == io_addr ? mem_367 : _GEN_1390; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1392 = 10'h170 == io_addr ? mem_368 : _GEN_1391; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1393 = 10'h171 == io_addr ? mem_369 : _GEN_1392; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1394 = 10'h172 == io_addr ? mem_370 : _GEN_1393; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1395 = 10'h173 == io_addr ? mem_371 : _GEN_1394; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1396 = 10'h174 == io_addr ? mem_372 : _GEN_1395; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1397 = 10'h175 == io_addr ? mem_373 : _GEN_1396; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1398 = 10'h176 == io_addr ? mem_374 : _GEN_1397; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1399 = 10'h177 == io_addr ? mem_375 : _GEN_1398; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1400 = 10'h178 == io_addr ? mem_376 : _GEN_1399; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1401 = 10'h179 == io_addr ? mem_377 : _GEN_1400; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1402 = 10'h17a == io_addr ? mem_378 : _GEN_1401; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1403 = 10'h17b == io_addr ? mem_379 : _GEN_1402; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1404 = 10'h17c == io_addr ? mem_380 : _GEN_1403; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1405 = 10'h17d == io_addr ? mem_381 : _GEN_1404; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1406 = 10'h17e == io_addr ? mem_382 : _GEN_1405; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1407 = 10'h17f == io_addr ? mem_383 : _GEN_1406; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1408 = 10'h180 == io_addr ? mem_384 : _GEN_1407; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1409 = 10'h181 == io_addr ? mem_385 : _GEN_1408; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1410 = 10'h182 == io_addr ? mem_386 : _GEN_1409; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1411 = 10'h183 == io_addr ? mem_387 : _GEN_1410; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1412 = 10'h184 == io_addr ? mem_388 : _GEN_1411; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1413 = 10'h185 == io_addr ? mem_389 : _GEN_1412; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1414 = 10'h186 == io_addr ? mem_390 : _GEN_1413; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1415 = 10'h187 == io_addr ? mem_391 : _GEN_1414; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1416 = 10'h188 == io_addr ? mem_392 : _GEN_1415; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1417 = 10'h189 == io_addr ? mem_393 : _GEN_1416; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1418 = 10'h18a == io_addr ? mem_394 : _GEN_1417; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1419 = 10'h18b == io_addr ? mem_395 : _GEN_1418; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1420 = 10'h18c == io_addr ? mem_396 : _GEN_1419; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1421 = 10'h18d == io_addr ? mem_397 : _GEN_1420; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1422 = 10'h18e == io_addr ? mem_398 : _GEN_1421; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1423 = 10'h18f == io_addr ? mem_399 : _GEN_1422; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1424 = 10'h190 == io_addr ? mem_400 : _GEN_1423; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1425 = 10'h191 == io_addr ? mem_401 : _GEN_1424; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1426 = 10'h192 == io_addr ? mem_402 : _GEN_1425; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1427 = 10'h193 == io_addr ? mem_403 : _GEN_1426; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1428 = 10'h194 == io_addr ? mem_404 : _GEN_1427; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1429 = 10'h195 == io_addr ? mem_405 : _GEN_1428; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1430 = 10'h196 == io_addr ? mem_406 : _GEN_1429; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1431 = 10'h197 == io_addr ? mem_407 : _GEN_1430; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1432 = 10'h198 == io_addr ? mem_408 : _GEN_1431; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1433 = 10'h199 == io_addr ? mem_409 : _GEN_1432; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1434 = 10'h19a == io_addr ? mem_410 : _GEN_1433; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1435 = 10'h19b == io_addr ? mem_411 : _GEN_1434; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1436 = 10'h19c == io_addr ? mem_412 : _GEN_1435; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1437 = 10'h19d == io_addr ? mem_413 : _GEN_1436; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1438 = 10'h19e == io_addr ? mem_414 : _GEN_1437; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1439 = 10'h19f == io_addr ? mem_415 : _GEN_1438; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1440 = 10'h1a0 == io_addr ? mem_416 : _GEN_1439; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1441 = 10'h1a1 == io_addr ? mem_417 : _GEN_1440; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1442 = 10'h1a2 == io_addr ? mem_418 : _GEN_1441; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1443 = 10'h1a3 == io_addr ? mem_419 : _GEN_1442; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1444 = 10'h1a4 == io_addr ? mem_420 : _GEN_1443; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1445 = 10'h1a5 == io_addr ? mem_421 : _GEN_1444; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1446 = 10'h1a6 == io_addr ? mem_422 : _GEN_1445; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1447 = 10'h1a7 == io_addr ? mem_423 : _GEN_1446; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1448 = 10'h1a8 == io_addr ? mem_424 : _GEN_1447; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1449 = 10'h1a9 == io_addr ? mem_425 : _GEN_1448; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1450 = 10'h1aa == io_addr ? mem_426 : _GEN_1449; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1451 = 10'h1ab == io_addr ? mem_427 : _GEN_1450; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1452 = 10'h1ac == io_addr ? mem_428 : _GEN_1451; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1453 = 10'h1ad == io_addr ? mem_429 : _GEN_1452; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1454 = 10'h1ae == io_addr ? mem_430 : _GEN_1453; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1455 = 10'h1af == io_addr ? mem_431 : _GEN_1454; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1456 = 10'h1b0 == io_addr ? mem_432 : _GEN_1455; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1457 = 10'h1b1 == io_addr ? mem_433 : _GEN_1456; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1458 = 10'h1b2 == io_addr ? mem_434 : _GEN_1457; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1459 = 10'h1b3 == io_addr ? mem_435 : _GEN_1458; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1460 = 10'h1b4 == io_addr ? mem_436 : _GEN_1459; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1461 = 10'h1b5 == io_addr ? mem_437 : _GEN_1460; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1462 = 10'h1b6 == io_addr ? mem_438 : _GEN_1461; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1463 = 10'h1b7 == io_addr ? mem_439 : _GEN_1462; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1464 = 10'h1b8 == io_addr ? mem_440 : _GEN_1463; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1465 = 10'h1b9 == io_addr ? mem_441 : _GEN_1464; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1466 = 10'h1ba == io_addr ? mem_442 : _GEN_1465; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1467 = 10'h1bb == io_addr ? mem_443 : _GEN_1466; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1468 = 10'h1bc == io_addr ? mem_444 : _GEN_1467; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1469 = 10'h1bd == io_addr ? mem_445 : _GEN_1468; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1470 = 10'h1be == io_addr ? mem_446 : _GEN_1469; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1471 = 10'h1bf == io_addr ? mem_447 : _GEN_1470; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1472 = 10'h1c0 == io_addr ? mem_448 : _GEN_1471; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1473 = 10'h1c1 == io_addr ? mem_449 : _GEN_1472; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1474 = 10'h1c2 == io_addr ? mem_450 : _GEN_1473; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1475 = 10'h1c3 == io_addr ? mem_451 : _GEN_1474; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1476 = 10'h1c4 == io_addr ? mem_452 : _GEN_1475; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1477 = 10'h1c5 == io_addr ? mem_453 : _GEN_1476; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1478 = 10'h1c6 == io_addr ? mem_454 : _GEN_1477; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1479 = 10'h1c7 == io_addr ? mem_455 : _GEN_1478; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1480 = 10'h1c8 == io_addr ? mem_456 : _GEN_1479; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1481 = 10'h1c9 == io_addr ? mem_457 : _GEN_1480; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1482 = 10'h1ca == io_addr ? mem_458 : _GEN_1481; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1483 = 10'h1cb == io_addr ? mem_459 : _GEN_1482; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1484 = 10'h1cc == io_addr ? mem_460 : _GEN_1483; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1485 = 10'h1cd == io_addr ? mem_461 : _GEN_1484; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1486 = 10'h1ce == io_addr ? mem_462 : _GEN_1485; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1487 = 10'h1cf == io_addr ? mem_463 : _GEN_1486; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1488 = 10'h1d0 == io_addr ? mem_464 : _GEN_1487; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1489 = 10'h1d1 == io_addr ? mem_465 : _GEN_1488; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1490 = 10'h1d2 == io_addr ? mem_466 : _GEN_1489; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1491 = 10'h1d3 == io_addr ? mem_467 : _GEN_1490; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1492 = 10'h1d4 == io_addr ? mem_468 : _GEN_1491; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1493 = 10'h1d5 == io_addr ? mem_469 : _GEN_1492; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1494 = 10'h1d6 == io_addr ? mem_470 : _GEN_1493; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1495 = 10'h1d7 == io_addr ? mem_471 : _GEN_1494; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1496 = 10'h1d8 == io_addr ? mem_472 : _GEN_1495; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1497 = 10'h1d9 == io_addr ? mem_473 : _GEN_1496; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1498 = 10'h1da == io_addr ? mem_474 : _GEN_1497; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1499 = 10'h1db == io_addr ? mem_475 : _GEN_1498; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1500 = 10'h1dc == io_addr ? mem_476 : _GEN_1499; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1501 = 10'h1dd == io_addr ? mem_477 : _GEN_1500; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1502 = 10'h1de == io_addr ? mem_478 : _GEN_1501; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1503 = 10'h1df == io_addr ? mem_479 : _GEN_1502; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1504 = 10'h1e0 == io_addr ? mem_480 : _GEN_1503; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1505 = 10'h1e1 == io_addr ? mem_481 : _GEN_1504; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1506 = 10'h1e2 == io_addr ? mem_482 : _GEN_1505; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1507 = 10'h1e3 == io_addr ? mem_483 : _GEN_1506; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1508 = 10'h1e4 == io_addr ? mem_484 : _GEN_1507; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1509 = 10'h1e5 == io_addr ? mem_485 : _GEN_1508; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1510 = 10'h1e6 == io_addr ? mem_486 : _GEN_1509; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1511 = 10'h1e7 == io_addr ? mem_487 : _GEN_1510; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1512 = 10'h1e8 == io_addr ? mem_488 : _GEN_1511; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1513 = 10'h1e9 == io_addr ? mem_489 : _GEN_1512; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1514 = 10'h1ea == io_addr ? mem_490 : _GEN_1513; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1515 = 10'h1eb == io_addr ? mem_491 : _GEN_1514; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1516 = 10'h1ec == io_addr ? mem_492 : _GEN_1515; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1517 = 10'h1ed == io_addr ? mem_493 : _GEN_1516; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1518 = 10'h1ee == io_addr ? mem_494 : _GEN_1517; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1519 = 10'h1ef == io_addr ? mem_495 : _GEN_1518; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1520 = 10'h1f0 == io_addr ? mem_496 : _GEN_1519; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1521 = 10'h1f1 == io_addr ? mem_497 : _GEN_1520; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1522 = 10'h1f2 == io_addr ? mem_498 : _GEN_1521; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1523 = 10'h1f3 == io_addr ? mem_499 : _GEN_1522; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1524 = 10'h1f4 == io_addr ? mem_500 : _GEN_1523; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1525 = 10'h1f5 == io_addr ? mem_501 : _GEN_1524; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1526 = 10'h1f6 == io_addr ? mem_502 : _GEN_1525; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1527 = 10'h1f7 == io_addr ? mem_503 : _GEN_1526; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1528 = 10'h1f8 == io_addr ? mem_504 : _GEN_1527; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1529 = 10'h1f9 == io_addr ? mem_505 : _GEN_1528; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1530 = 10'h1fa == io_addr ? mem_506 : _GEN_1529; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1531 = 10'h1fb == io_addr ? mem_507 : _GEN_1530; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1532 = 10'h1fc == io_addr ? mem_508 : _GEN_1531; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1533 = 10'h1fd == io_addr ? mem_509 : _GEN_1532; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1534 = 10'h1fe == io_addr ? mem_510 : _GEN_1533; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1535 = 10'h1ff == io_addr ? mem_511 : _GEN_1534; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1536 = 10'h200 == io_addr ? mem_512 : _GEN_1535; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1537 = 10'h201 == io_addr ? mem_513 : _GEN_1536; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1538 = 10'h202 == io_addr ? mem_514 : _GEN_1537; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1539 = 10'h203 == io_addr ? mem_515 : _GEN_1538; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1540 = 10'h204 == io_addr ? mem_516 : _GEN_1539; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1541 = 10'h205 == io_addr ? mem_517 : _GEN_1540; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1542 = 10'h206 == io_addr ? mem_518 : _GEN_1541; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1543 = 10'h207 == io_addr ? mem_519 : _GEN_1542; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1544 = 10'h208 == io_addr ? mem_520 : _GEN_1543; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1545 = 10'h209 == io_addr ? mem_521 : _GEN_1544; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1546 = 10'h20a == io_addr ? mem_522 : _GEN_1545; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1547 = 10'h20b == io_addr ? mem_523 : _GEN_1546; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1548 = 10'h20c == io_addr ? mem_524 : _GEN_1547; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1549 = 10'h20d == io_addr ? mem_525 : _GEN_1548; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1550 = 10'h20e == io_addr ? mem_526 : _GEN_1549; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1551 = 10'h20f == io_addr ? mem_527 : _GEN_1550; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1552 = 10'h210 == io_addr ? mem_528 : _GEN_1551; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1553 = 10'h211 == io_addr ? mem_529 : _GEN_1552; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1554 = 10'h212 == io_addr ? mem_530 : _GEN_1553; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1555 = 10'h213 == io_addr ? mem_531 : _GEN_1554; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1556 = 10'h214 == io_addr ? mem_532 : _GEN_1555; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1557 = 10'h215 == io_addr ? mem_533 : _GEN_1556; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1558 = 10'h216 == io_addr ? mem_534 : _GEN_1557; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1559 = 10'h217 == io_addr ? mem_535 : _GEN_1558; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1560 = 10'h218 == io_addr ? mem_536 : _GEN_1559; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1561 = 10'h219 == io_addr ? mem_537 : _GEN_1560; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1562 = 10'h21a == io_addr ? mem_538 : _GEN_1561; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1563 = 10'h21b == io_addr ? mem_539 : _GEN_1562; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1564 = 10'h21c == io_addr ? mem_540 : _GEN_1563; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1565 = 10'h21d == io_addr ? mem_541 : _GEN_1564; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1566 = 10'h21e == io_addr ? mem_542 : _GEN_1565; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1567 = 10'h21f == io_addr ? mem_543 : _GEN_1566; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1568 = 10'h220 == io_addr ? mem_544 : _GEN_1567; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1569 = 10'h221 == io_addr ? mem_545 : _GEN_1568; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1570 = 10'h222 == io_addr ? mem_546 : _GEN_1569; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1571 = 10'h223 == io_addr ? mem_547 : _GEN_1570; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1572 = 10'h224 == io_addr ? mem_548 : _GEN_1571; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1573 = 10'h225 == io_addr ? mem_549 : _GEN_1572; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1574 = 10'h226 == io_addr ? mem_550 : _GEN_1573; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1575 = 10'h227 == io_addr ? mem_551 : _GEN_1574; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1576 = 10'h228 == io_addr ? mem_552 : _GEN_1575; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1577 = 10'h229 == io_addr ? mem_553 : _GEN_1576; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1578 = 10'h22a == io_addr ? mem_554 : _GEN_1577; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1579 = 10'h22b == io_addr ? mem_555 : _GEN_1578; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1580 = 10'h22c == io_addr ? mem_556 : _GEN_1579; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1581 = 10'h22d == io_addr ? mem_557 : _GEN_1580; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1582 = 10'h22e == io_addr ? mem_558 : _GEN_1581; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1583 = 10'h22f == io_addr ? mem_559 : _GEN_1582; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1584 = 10'h230 == io_addr ? mem_560 : _GEN_1583; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1585 = 10'h231 == io_addr ? mem_561 : _GEN_1584; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1586 = 10'h232 == io_addr ? mem_562 : _GEN_1585; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1587 = 10'h233 == io_addr ? mem_563 : _GEN_1586; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1588 = 10'h234 == io_addr ? mem_564 : _GEN_1587; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1589 = 10'h235 == io_addr ? mem_565 : _GEN_1588; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1590 = 10'h236 == io_addr ? mem_566 : _GEN_1589; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1591 = 10'h237 == io_addr ? mem_567 : _GEN_1590; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1592 = 10'h238 == io_addr ? mem_568 : _GEN_1591; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1593 = 10'h239 == io_addr ? mem_569 : _GEN_1592; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1594 = 10'h23a == io_addr ? mem_570 : _GEN_1593; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1595 = 10'h23b == io_addr ? mem_571 : _GEN_1594; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1596 = 10'h23c == io_addr ? mem_572 : _GEN_1595; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1597 = 10'h23d == io_addr ? mem_573 : _GEN_1596; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1598 = 10'h23e == io_addr ? mem_574 : _GEN_1597; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1599 = 10'h23f == io_addr ? mem_575 : _GEN_1598; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1600 = 10'h240 == io_addr ? mem_576 : _GEN_1599; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1601 = 10'h241 == io_addr ? mem_577 : _GEN_1600; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1602 = 10'h242 == io_addr ? mem_578 : _GEN_1601; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1603 = 10'h243 == io_addr ? mem_579 : _GEN_1602; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1604 = 10'h244 == io_addr ? mem_580 : _GEN_1603; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1605 = 10'h245 == io_addr ? mem_581 : _GEN_1604; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1606 = 10'h246 == io_addr ? mem_582 : _GEN_1605; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1607 = 10'h247 == io_addr ? mem_583 : _GEN_1606; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1608 = 10'h248 == io_addr ? mem_584 : _GEN_1607; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1609 = 10'h249 == io_addr ? mem_585 : _GEN_1608; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1610 = 10'h24a == io_addr ? mem_586 : _GEN_1609; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1611 = 10'h24b == io_addr ? mem_587 : _GEN_1610; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1612 = 10'h24c == io_addr ? mem_588 : _GEN_1611; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1613 = 10'h24d == io_addr ? mem_589 : _GEN_1612; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1614 = 10'h24e == io_addr ? mem_590 : _GEN_1613; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1615 = 10'h24f == io_addr ? mem_591 : _GEN_1614; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1616 = 10'h250 == io_addr ? mem_592 : _GEN_1615; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1617 = 10'h251 == io_addr ? mem_593 : _GEN_1616; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1618 = 10'h252 == io_addr ? mem_594 : _GEN_1617; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1619 = 10'h253 == io_addr ? mem_595 : _GEN_1618; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1620 = 10'h254 == io_addr ? mem_596 : _GEN_1619; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1621 = 10'h255 == io_addr ? mem_597 : _GEN_1620; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1622 = 10'h256 == io_addr ? mem_598 : _GEN_1621; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1623 = 10'h257 == io_addr ? mem_599 : _GEN_1622; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1624 = 10'h258 == io_addr ? mem_600 : _GEN_1623; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1625 = 10'h259 == io_addr ? mem_601 : _GEN_1624; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1626 = 10'h25a == io_addr ? mem_602 : _GEN_1625; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1627 = 10'h25b == io_addr ? mem_603 : _GEN_1626; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1628 = 10'h25c == io_addr ? mem_604 : _GEN_1627; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1629 = 10'h25d == io_addr ? mem_605 : _GEN_1628; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1630 = 10'h25e == io_addr ? mem_606 : _GEN_1629; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1631 = 10'h25f == io_addr ? mem_607 : _GEN_1630; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1632 = 10'h260 == io_addr ? mem_608 : _GEN_1631; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1633 = 10'h261 == io_addr ? mem_609 : _GEN_1632; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1634 = 10'h262 == io_addr ? mem_610 : _GEN_1633; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1635 = 10'h263 == io_addr ? mem_611 : _GEN_1634; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1636 = 10'h264 == io_addr ? mem_612 : _GEN_1635; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1637 = 10'h265 == io_addr ? mem_613 : _GEN_1636; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1638 = 10'h266 == io_addr ? mem_614 : _GEN_1637; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1639 = 10'h267 == io_addr ? mem_615 : _GEN_1638; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1640 = 10'h268 == io_addr ? mem_616 : _GEN_1639; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1641 = 10'h269 == io_addr ? mem_617 : _GEN_1640; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1642 = 10'h26a == io_addr ? mem_618 : _GEN_1641; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1643 = 10'h26b == io_addr ? mem_619 : _GEN_1642; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1644 = 10'h26c == io_addr ? mem_620 : _GEN_1643; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1645 = 10'h26d == io_addr ? mem_621 : _GEN_1644; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1646 = 10'h26e == io_addr ? mem_622 : _GEN_1645; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1647 = 10'h26f == io_addr ? mem_623 : _GEN_1646; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1648 = 10'h270 == io_addr ? mem_624 : _GEN_1647; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1649 = 10'h271 == io_addr ? mem_625 : _GEN_1648; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1650 = 10'h272 == io_addr ? mem_626 : _GEN_1649; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1651 = 10'h273 == io_addr ? mem_627 : _GEN_1650; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1652 = 10'h274 == io_addr ? mem_628 : _GEN_1651; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1653 = 10'h275 == io_addr ? mem_629 : _GEN_1652; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1654 = 10'h276 == io_addr ? mem_630 : _GEN_1653; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1655 = 10'h277 == io_addr ? mem_631 : _GEN_1654; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1656 = 10'h278 == io_addr ? mem_632 : _GEN_1655; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1657 = 10'h279 == io_addr ? mem_633 : _GEN_1656; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1658 = 10'h27a == io_addr ? mem_634 : _GEN_1657; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1659 = 10'h27b == io_addr ? mem_635 : _GEN_1658; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1660 = 10'h27c == io_addr ? mem_636 : _GEN_1659; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1661 = 10'h27d == io_addr ? mem_637 : _GEN_1660; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1662 = 10'h27e == io_addr ? mem_638 : _GEN_1661; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1663 = 10'h27f == io_addr ? mem_639 : _GEN_1662; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1664 = 10'h280 == io_addr ? mem_640 : _GEN_1663; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1665 = 10'h281 == io_addr ? mem_641 : _GEN_1664; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1666 = 10'h282 == io_addr ? mem_642 : _GEN_1665; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1667 = 10'h283 == io_addr ? mem_643 : _GEN_1666; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1668 = 10'h284 == io_addr ? mem_644 : _GEN_1667; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1669 = 10'h285 == io_addr ? mem_645 : _GEN_1668; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1670 = 10'h286 == io_addr ? mem_646 : _GEN_1669; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1671 = 10'h287 == io_addr ? mem_647 : _GEN_1670; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1672 = 10'h288 == io_addr ? mem_648 : _GEN_1671; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1673 = 10'h289 == io_addr ? mem_649 : _GEN_1672; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1674 = 10'h28a == io_addr ? mem_650 : _GEN_1673; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1675 = 10'h28b == io_addr ? mem_651 : _GEN_1674; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1676 = 10'h28c == io_addr ? mem_652 : _GEN_1675; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1677 = 10'h28d == io_addr ? mem_653 : _GEN_1676; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1678 = 10'h28e == io_addr ? mem_654 : _GEN_1677; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1679 = 10'h28f == io_addr ? mem_655 : _GEN_1678; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1680 = 10'h290 == io_addr ? mem_656 : _GEN_1679; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1681 = 10'h291 == io_addr ? mem_657 : _GEN_1680; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1682 = 10'h292 == io_addr ? mem_658 : _GEN_1681; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1683 = 10'h293 == io_addr ? mem_659 : _GEN_1682; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1684 = 10'h294 == io_addr ? mem_660 : _GEN_1683; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1685 = 10'h295 == io_addr ? mem_661 : _GEN_1684; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1686 = 10'h296 == io_addr ? mem_662 : _GEN_1685; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1687 = 10'h297 == io_addr ? mem_663 : _GEN_1686; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1688 = 10'h298 == io_addr ? mem_664 : _GEN_1687; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1689 = 10'h299 == io_addr ? mem_665 : _GEN_1688; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1690 = 10'h29a == io_addr ? mem_666 : _GEN_1689; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1691 = 10'h29b == io_addr ? mem_667 : _GEN_1690; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1692 = 10'h29c == io_addr ? mem_668 : _GEN_1691; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1693 = 10'h29d == io_addr ? mem_669 : _GEN_1692; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1694 = 10'h29e == io_addr ? mem_670 : _GEN_1693; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1695 = 10'h29f == io_addr ? mem_671 : _GEN_1694; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1696 = 10'h2a0 == io_addr ? mem_672 : _GEN_1695; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1697 = 10'h2a1 == io_addr ? mem_673 : _GEN_1696; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1698 = 10'h2a2 == io_addr ? mem_674 : _GEN_1697; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1699 = 10'h2a3 == io_addr ? mem_675 : _GEN_1698; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1700 = 10'h2a4 == io_addr ? mem_676 : _GEN_1699; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1701 = 10'h2a5 == io_addr ? mem_677 : _GEN_1700; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1702 = 10'h2a6 == io_addr ? mem_678 : _GEN_1701; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1703 = 10'h2a7 == io_addr ? mem_679 : _GEN_1702; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1704 = 10'h2a8 == io_addr ? mem_680 : _GEN_1703; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1705 = 10'h2a9 == io_addr ? mem_681 : _GEN_1704; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1706 = 10'h2aa == io_addr ? mem_682 : _GEN_1705; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1707 = 10'h2ab == io_addr ? mem_683 : _GEN_1706; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1708 = 10'h2ac == io_addr ? mem_684 : _GEN_1707; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1709 = 10'h2ad == io_addr ? mem_685 : _GEN_1708; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1710 = 10'h2ae == io_addr ? mem_686 : _GEN_1709; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1711 = 10'h2af == io_addr ? mem_687 : _GEN_1710; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1712 = 10'h2b0 == io_addr ? mem_688 : _GEN_1711; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1713 = 10'h2b1 == io_addr ? mem_689 : _GEN_1712; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1714 = 10'h2b2 == io_addr ? mem_690 : _GEN_1713; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1715 = 10'h2b3 == io_addr ? mem_691 : _GEN_1714; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1716 = 10'h2b4 == io_addr ? mem_692 : _GEN_1715; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1717 = 10'h2b5 == io_addr ? mem_693 : _GEN_1716; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1718 = 10'h2b6 == io_addr ? mem_694 : _GEN_1717; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1719 = 10'h2b7 == io_addr ? mem_695 : _GEN_1718; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1720 = 10'h2b8 == io_addr ? mem_696 : _GEN_1719; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1721 = 10'h2b9 == io_addr ? mem_697 : _GEN_1720; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1722 = 10'h2ba == io_addr ? mem_698 : _GEN_1721; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1723 = 10'h2bb == io_addr ? mem_699 : _GEN_1722; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1724 = 10'h2bc == io_addr ? mem_700 : _GEN_1723; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1725 = 10'h2bd == io_addr ? mem_701 : _GEN_1724; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1726 = 10'h2be == io_addr ? mem_702 : _GEN_1725; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1727 = 10'h2bf == io_addr ? mem_703 : _GEN_1726; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1728 = 10'h2c0 == io_addr ? mem_704 : _GEN_1727; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1729 = 10'h2c1 == io_addr ? mem_705 : _GEN_1728; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1730 = 10'h2c2 == io_addr ? mem_706 : _GEN_1729; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1731 = 10'h2c3 == io_addr ? mem_707 : _GEN_1730; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1732 = 10'h2c4 == io_addr ? mem_708 : _GEN_1731; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1733 = 10'h2c5 == io_addr ? mem_709 : _GEN_1732; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1734 = 10'h2c6 == io_addr ? mem_710 : _GEN_1733; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1735 = 10'h2c7 == io_addr ? mem_711 : _GEN_1734; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1736 = 10'h2c8 == io_addr ? mem_712 : _GEN_1735; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1737 = 10'h2c9 == io_addr ? mem_713 : _GEN_1736; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1738 = 10'h2ca == io_addr ? mem_714 : _GEN_1737; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1739 = 10'h2cb == io_addr ? mem_715 : _GEN_1738; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1740 = 10'h2cc == io_addr ? mem_716 : _GEN_1739; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1741 = 10'h2cd == io_addr ? mem_717 : _GEN_1740; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1742 = 10'h2ce == io_addr ? mem_718 : _GEN_1741; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1743 = 10'h2cf == io_addr ? mem_719 : _GEN_1742; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1744 = 10'h2d0 == io_addr ? mem_720 : _GEN_1743; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1745 = 10'h2d1 == io_addr ? mem_721 : _GEN_1744; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1746 = 10'h2d2 == io_addr ? mem_722 : _GEN_1745; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1747 = 10'h2d3 == io_addr ? mem_723 : _GEN_1746; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1748 = 10'h2d4 == io_addr ? mem_724 : _GEN_1747; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1749 = 10'h2d5 == io_addr ? mem_725 : _GEN_1748; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1750 = 10'h2d6 == io_addr ? mem_726 : _GEN_1749; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1751 = 10'h2d7 == io_addr ? mem_727 : _GEN_1750; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1752 = 10'h2d8 == io_addr ? mem_728 : _GEN_1751; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1753 = 10'h2d9 == io_addr ? mem_729 : _GEN_1752; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1754 = 10'h2da == io_addr ? mem_730 : _GEN_1753; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1755 = 10'h2db == io_addr ? mem_731 : _GEN_1754; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1756 = 10'h2dc == io_addr ? mem_732 : _GEN_1755; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1757 = 10'h2dd == io_addr ? mem_733 : _GEN_1756; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1758 = 10'h2de == io_addr ? mem_734 : _GEN_1757; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1759 = 10'h2df == io_addr ? mem_735 : _GEN_1758; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1760 = 10'h2e0 == io_addr ? mem_736 : _GEN_1759; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1761 = 10'h2e1 == io_addr ? mem_737 : _GEN_1760; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1762 = 10'h2e2 == io_addr ? mem_738 : _GEN_1761; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1763 = 10'h2e3 == io_addr ? mem_739 : _GEN_1762; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1764 = 10'h2e4 == io_addr ? mem_740 : _GEN_1763; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1765 = 10'h2e5 == io_addr ? mem_741 : _GEN_1764; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1766 = 10'h2e6 == io_addr ? mem_742 : _GEN_1765; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1767 = 10'h2e7 == io_addr ? mem_743 : _GEN_1766; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1768 = 10'h2e8 == io_addr ? mem_744 : _GEN_1767; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1769 = 10'h2e9 == io_addr ? mem_745 : _GEN_1768; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1770 = 10'h2ea == io_addr ? mem_746 : _GEN_1769; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1771 = 10'h2eb == io_addr ? mem_747 : _GEN_1770; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1772 = 10'h2ec == io_addr ? mem_748 : _GEN_1771; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1773 = 10'h2ed == io_addr ? mem_749 : _GEN_1772; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1774 = 10'h2ee == io_addr ? mem_750 : _GEN_1773; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1775 = 10'h2ef == io_addr ? mem_751 : _GEN_1774; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1776 = 10'h2f0 == io_addr ? mem_752 : _GEN_1775; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1777 = 10'h2f1 == io_addr ? mem_753 : _GEN_1776; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1778 = 10'h2f2 == io_addr ? mem_754 : _GEN_1777; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1779 = 10'h2f3 == io_addr ? mem_755 : _GEN_1778; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1780 = 10'h2f4 == io_addr ? mem_756 : _GEN_1779; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1781 = 10'h2f5 == io_addr ? mem_757 : _GEN_1780; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1782 = 10'h2f6 == io_addr ? mem_758 : _GEN_1781; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1783 = 10'h2f7 == io_addr ? mem_759 : _GEN_1782; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1784 = 10'h2f8 == io_addr ? mem_760 : _GEN_1783; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1785 = 10'h2f9 == io_addr ? mem_761 : _GEN_1784; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1786 = 10'h2fa == io_addr ? mem_762 : _GEN_1785; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1787 = 10'h2fb == io_addr ? mem_763 : _GEN_1786; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1788 = 10'h2fc == io_addr ? mem_764 : _GEN_1787; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1789 = 10'h2fd == io_addr ? mem_765 : _GEN_1788; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1790 = 10'h2fe == io_addr ? mem_766 : _GEN_1789; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1791 = 10'h2ff == io_addr ? mem_767 : _GEN_1790; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1792 = 10'h300 == io_addr ? mem_768 : _GEN_1791; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1793 = 10'h301 == io_addr ? mem_769 : _GEN_1792; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1794 = 10'h302 == io_addr ? mem_770 : _GEN_1793; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1795 = 10'h303 == io_addr ? mem_771 : _GEN_1794; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1796 = 10'h304 == io_addr ? mem_772 : _GEN_1795; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1797 = 10'h305 == io_addr ? mem_773 : _GEN_1796; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1798 = 10'h306 == io_addr ? mem_774 : _GEN_1797; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1799 = 10'h307 == io_addr ? mem_775 : _GEN_1798; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1800 = 10'h308 == io_addr ? mem_776 : _GEN_1799; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1801 = 10'h309 == io_addr ? mem_777 : _GEN_1800; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1802 = 10'h30a == io_addr ? mem_778 : _GEN_1801; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1803 = 10'h30b == io_addr ? mem_779 : _GEN_1802; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1804 = 10'h30c == io_addr ? mem_780 : _GEN_1803; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1805 = 10'h30d == io_addr ? mem_781 : _GEN_1804; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1806 = 10'h30e == io_addr ? mem_782 : _GEN_1805; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1807 = 10'h30f == io_addr ? mem_783 : _GEN_1806; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1808 = 10'h310 == io_addr ? mem_784 : _GEN_1807; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1809 = 10'h311 == io_addr ? mem_785 : _GEN_1808; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1810 = 10'h312 == io_addr ? mem_786 : _GEN_1809; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1811 = 10'h313 == io_addr ? mem_787 : _GEN_1810; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1812 = 10'h314 == io_addr ? mem_788 : _GEN_1811; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1813 = 10'h315 == io_addr ? mem_789 : _GEN_1812; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1814 = 10'h316 == io_addr ? mem_790 : _GEN_1813; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1815 = 10'h317 == io_addr ? mem_791 : _GEN_1814; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1816 = 10'h318 == io_addr ? mem_792 : _GEN_1815; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1817 = 10'h319 == io_addr ? mem_793 : _GEN_1816; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1818 = 10'h31a == io_addr ? mem_794 : _GEN_1817; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1819 = 10'h31b == io_addr ? mem_795 : _GEN_1818; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1820 = 10'h31c == io_addr ? mem_796 : _GEN_1819; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1821 = 10'h31d == io_addr ? mem_797 : _GEN_1820; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1822 = 10'h31e == io_addr ? mem_798 : _GEN_1821; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1823 = 10'h31f == io_addr ? mem_799 : _GEN_1822; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1824 = 10'h320 == io_addr ? mem_800 : _GEN_1823; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1825 = 10'h321 == io_addr ? mem_801 : _GEN_1824; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1826 = 10'h322 == io_addr ? mem_802 : _GEN_1825; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1827 = 10'h323 == io_addr ? mem_803 : _GEN_1826; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1828 = 10'h324 == io_addr ? mem_804 : _GEN_1827; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1829 = 10'h325 == io_addr ? mem_805 : _GEN_1828; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1830 = 10'h326 == io_addr ? mem_806 : _GEN_1829; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1831 = 10'h327 == io_addr ? mem_807 : _GEN_1830; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1832 = 10'h328 == io_addr ? mem_808 : _GEN_1831; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1833 = 10'h329 == io_addr ? mem_809 : _GEN_1832; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1834 = 10'h32a == io_addr ? mem_810 : _GEN_1833; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1835 = 10'h32b == io_addr ? mem_811 : _GEN_1834; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1836 = 10'h32c == io_addr ? mem_812 : _GEN_1835; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1837 = 10'h32d == io_addr ? mem_813 : _GEN_1836; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1838 = 10'h32e == io_addr ? mem_814 : _GEN_1837; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1839 = 10'h32f == io_addr ? mem_815 : _GEN_1838; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1840 = 10'h330 == io_addr ? mem_816 : _GEN_1839; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1841 = 10'h331 == io_addr ? mem_817 : _GEN_1840; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1842 = 10'h332 == io_addr ? mem_818 : _GEN_1841; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1843 = 10'h333 == io_addr ? mem_819 : _GEN_1842; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1844 = 10'h334 == io_addr ? mem_820 : _GEN_1843; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1845 = 10'h335 == io_addr ? mem_821 : _GEN_1844; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1846 = 10'h336 == io_addr ? mem_822 : _GEN_1845; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1847 = 10'h337 == io_addr ? mem_823 : _GEN_1846; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1848 = 10'h338 == io_addr ? mem_824 : _GEN_1847; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1849 = 10'h339 == io_addr ? mem_825 : _GEN_1848; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1850 = 10'h33a == io_addr ? mem_826 : _GEN_1849; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1851 = 10'h33b == io_addr ? mem_827 : _GEN_1850; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1852 = 10'h33c == io_addr ? mem_828 : _GEN_1851; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1853 = 10'h33d == io_addr ? mem_829 : _GEN_1852; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1854 = 10'h33e == io_addr ? mem_830 : _GEN_1853; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1855 = 10'h33f == io_addr ? mem_831 : _GEN_1854; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1856 = 10'h340 == io_addr ? mem_832 : _GEN_1855; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1857 = 10'h341 == io_addr ? mem_833 : _GEN_1856; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1858 = 10'h342 == io_addr ? mem_834 : _GEN_1857; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1859 = 10'h343 == io_addr ? mem_835 : _GEN_1858; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1860 = 10'h344 == io_addr ? mem_836 : _GEN_1859; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1861 = 10'h345 == io_addr ? mem_837 : _GEN_1860; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1862 = 10'h346 == io_addr ? mem_838 : _GEN_1861; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1863 = 10'h347 == io_addr ? mem_839 : _GEN_1862; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1864 = 10'h348 == io_addr ? mem_840 : _GEN_1863; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1865 = 10'h349 == io_addr ? mem_841 : _GEN_1864; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1866 = 10'h34a == io_addr ? mem_842 : _GEN_1865; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1867 = 10'h34b == io_addr ? mem_843 : _GEN_1866; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1868 = 10'h34c == io_addr ? mem_844 : _GEN_1867; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1869 = 10'h34d == io_addr ? mem_845 : _GEN_1868; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1870 = 10'h34e == io_addr ? mem_846 : _GEN_1869; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1871 = 10'h34f == io_addr ? mem_847 : _GEN_1870; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1872 = 10'h350 == io_addr ? mem_848 : _GEN_1871; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1873 = 10'h351 == io_addr ? mem_849 : _GEN_1872; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1874 = 10'h352 == io_addr ? mem_850 : _GEN_1873; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1875 = 10'h353 == io_addr ? mem_851 : _GEN_1874; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1876 = 10'h354 == io_addr ? mem_852 : _GEN_1875; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1877 = 10'h355 == io_addr ? mem_853 : _GEN_1876; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1878 = 10'h356 == io_addr ? mem_854 : _GEN_1877; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1879 = 10'h357 == io_addr ? mem_855 : _GEN_1878; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1880 = 10'h358 == io_addr ? mem_856 : _GEN_1879; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1881 = 10'h359 == io_addr ? mem_857 : _GEN_1880; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1882 = 10'h35a == io_addr ? mem_858 : _GEN_1881; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1883 = 10'h35b == io_addr ? mem_859 : _GEN_1882; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1884 = 10'h35c == io_addr ? mem_860 : _GEN_1883; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1885 = 10'h35d == io_addr ? mem_861 : _GEN_1884; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1886 = 10'h35e == io_addr ? mem_862 : _GEN_1885; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1887 = 10'h35f == io_addr ? mem_863 : _GEN_1886; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1888 = 10'h360 == io_addr ? mem_864 : _GEN_1887; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1889 = 10'h361 == io_addr ? mem_865 : _GEN_1888; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1890 = 10'h362 == io_addr ? mem_866 : _GEN_1889; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1891 = 10'h363 == io_addr ? mem_867 : _GEN_1890; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1892 = 10'h364 == io_addr ? mem_868 : _GEN_1891; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1893 = 10'h365 == io_addr ? mem_869 : _GEN_1892; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1894 = 10'h366 == io_addr ? mem_870 : _GEN_1893; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1895 = 10'h367 == io_addr ? mem_871 : _GEN_1894; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1896 = 10'h368 == io_addr ? mem_872 : _GEN_1895; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1897 = 10'h369 == io_addr ? mem_873 : _GEN_1896; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1898 = 10'h36a == io_addr ? mem_874 : _GEN_1897; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1899 = 10'h36b == io_addr ? mem_875 : _GEN_1898; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1900 = 10'h36c == io_addr ? mem_876 : _GEN_1899; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1901 = 10'h36d == io_addr ? mem_877 : _GEN_1900; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1902 = 10'h36e == io_addr ? mem_878 : _GEN_1901; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1903 = 10'h36f == io_addr ? mem_879 : _GEN_1902; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1904 = 10'h370 == io_addr ? mem_880 : _GEN_1903; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1905 = 10'h371 == io_addr ? mem_881 : _GEN_1904; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1906 = 10'h372 == io_addr ? mem_882 : _GEN_1905; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1907 = 10'h373 == io_addr ? mem_883 : _GEN_1906; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1908 = 10'h374 == io_addr ? mem_884 : _GEN_1907; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1909 = 10'h375 == io_addr ? mem_885 : _GEN_1908; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1910 = 10'h376 == io_addr ? mem_886 : _GEN_1909; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1911 = 10'h377 == io_addr ? mem_887 : _GEN_1910; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1912 = 10'h378 == io_addr ? mem_888 : _GEN_1911; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1913 = 10'h379 == io_addr ? mem_889 : _GEN_1912; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1914 = 10'h37a == io_addr ? mem_890 : _GEN_1913; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1915 = 10'h37b == io_addr ? mem_891 : _GEN_1914; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1916 = 10'h37c == io_addr ? mem_892 : _GEN_1915; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1917 = 10'h37d == io_addr ? mem_893 : _GEN_1916; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1918 = 10'h37e == io_addr ? mem_894 : _GEN_1917; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1919 = 10'h37f == io_addr ? mem_895 : _GEN_1918; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1920 = 10'h380 == io_addr ? mem_896 : _GEN_1919; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1921 = 10'h381 == io_addr ? mem_897 : _GEN_1920; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1922 = 10'h382 == io_addr ? mem_898 : _GEN_1921; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1923 = 10'h383 == io_addr ? mem_899 : _GEN_1922; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1924 = 10'h384 == io_addr ? mem_900 : _GEN_1923; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1925 = 10'h385 == io_addr ? mem_901 : _GEN_1924; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1926 = 10'h386 == io_addr ? mem_902 : _GEN_1925; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1927 = 10'h387 == io_addr ? mem_903 : _GEN_1926; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1928 = 10'h388 == io_addr ? mem_904 : _GEN_1927; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1929 = 10'h389 == io_addr ? mem_905 : _GEN_1928; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1930 = 10'h38a == io_addr ? mem_906 : _GEN_1929; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1931 = 10'h38b == io_addr ? mem_907 : _GEN_1930; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1932 = 10'h38c == io_addr ? mem_908 : _GEN_1931; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1933 = 10'h38d == io_addr ? mem_909 : _GEN_1932; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1934 = 10'h38e == io_addr ? mem_910 : _GEN_1933; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1935 = 10'h38f == io_addr ? mem_911 : _GEN_1934; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1936 = 10'h390 == io_addr ? mem_912 : _GEN_1935; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1937 = 10'h391 == io_addr ? mem_913 : _GEN_1936; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1938 = 10'h392 == io_addr ? mem_914 : _GEN_1937; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1939 = 10'h393 == io_addr ? mem_915 : _GEN_1938; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1940 = 10'h394 == io_addr ? mem_916 : _GEN_1939; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1941 = 10'h395 == io_addr ? mem_917 : _GEN_1940; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1942 = 10'h396 == io_addr ? mem_918 : _GEN_1941; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1943 = 10'h397 == io_addr ? mem_919 : _GEN_1942; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1944 = 10'h398 == io_addr ? mem_920 : _GEN_1943; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1945 = 10'h399 == io_addr ? mem_921 : _GEN_1944; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1946 = 10'h39a == io_addr ? mem_922 : _GEN_1945; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1947 = 10'h39b == io_addr ? mem_923 : _GEN_1946; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1948 = 10'h39c == io_addr ? mem_924 : _GEN_1947; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1949 = 10'h39d == io_addr ? mem_925 : _GEN_1948; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1950 = 10'h39e == io_addr ? mem_926 : _GEN_1949; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1951 = 10'h39f == io_addr ? mem_927 : _GEN_1950; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1952 = 10'h3a0 == io_addr ? mem_928 : _GEN_1951; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1953 = 10'h3a1 == io_addr ? mem_929 : _GEN_1952; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1954 = 10'h3a2 == io_addr ? mem_930 : _GEN_1953; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1955 = 10'h3a3 == io_addr ? mem_931 : _GEN_1954; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1956 = 10'h3a4 == io_addr ? mem_932 : _GEN_1955; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1957 = 10'h3a5 == io_addr ? mem_933 : _GEN_1956; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1958 = 10'h3a6 == io_addr ? mem_934 : _GEN_1957; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1959 = 10'h3a7 == io_addr ? mem_935 : _GEN_1958; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1960 = 10'h3a8 == io_addr ? mem_936 : _GEN_1959; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1961 = 10'h3a9 == io_addr ? mem_937 : _GEN_1960; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1962 = 10'h3aa == io_addr ? mem_938 : _GEN_1961; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1963 = 10'h3ab == io_addr ? mem_939 : _GEN_1962; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1964 = 10'h3ac == io_addr ? mem_940 : _GEN_1963; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1965 = 10'h3ad == io_addr ? mem_941 : _GEN_1964; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1966 = 10'h3ae == io_addr ? mem_942 : _GEN_1965; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1967 = 10'h3af == io_addr ? mem_943 : _GEN_1966; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1968 = 10'h3b0 == io_addr ? mem_944 : _GEN_1967; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1969 = 10'h3b1 == io_addr ? mem_945 : _GEN_1968; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1970 = 10'h3b2 == io_addr ? mem_946 : _GEN_1969; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1971 = 10'h3b3 == io_addr ? mem_947 : _GEN_1970; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1972 = 10'h3b4 == io_addr ? mem_948 : _GEN_1971; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1973 = 10'h3b5 == io_addr ? mem_949 : _GEN_1972; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1974 = 10'h3b6 == io_addr ? mem_950 : _GEN_1973; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1975 = 10'h3b7 == io_addr ? mem_951 : _GEN_1974; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1976 = 10'h3b8 == io_addr ? mem_952 : _GEN_1975; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1977 = 10'h3b9 == io_addr ? mem_953 : _GEN_1976; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1978 = 10'h3ba == io_addr ? mem_954 : _GEN_1977; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1979 = 10'h3bb == io_addr ? mem_955 : _GEN_1978; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1980 = 10'h3bc == io_addr ? mem_956 : _GEN_1979; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1981 = 10'h3bd == io_addr ? mem_957 : _GEN_1980; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1982 = 10'h3be == io_addr ? mem_958 : _GEN_1981; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1983 = 10'h3bf == io_addr ? mem_959 : _GEN_1982; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1984 = 10'h3c0 == io_addr ? mem_960 : _GEN_1983; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1985 = 10'h3c1 == io_addr ? mem_961 : _GEN_1984; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1986 = 10'h3c2 == io_addr ? mem_962 : _GEN_1985; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1987 = 10'h3c3 == io_addr ? mem_963 : _GEN_1986; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1988 = 10'h3c4 == io_addr ? mem_964 : _GEN_1987; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1989 = 10'h3c5 == io_addr ? mem_965 : _GEN_1988; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1990 = 10'h3c6 == io_addr ? mem_966 : _GEN_1989; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1991 = 10'h3c7 == io_addr ? mem_967 : _GEN_1990; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1992 = 10'h3c8 == io_addr ? mem_968 : _GEN_1991; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1993 = 10'h3c9 == io_addr ? mem_969 : _GEN_1992; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1994 = 10'h3ca == io_addr ? mem_970 : _GEN_1993; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1995 = 10'h3cb == io_addr ? mem_971 : _GEN_1994; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1996 = 10'h3cc == io_addr ? mem_972 : _GEN_1995; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1997 = 10'h3cd == io_addr ? mem_973 : _GEN_1996; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1998 = 10'h3ce == io_addr ? mem_974 : _GEN_1997; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_1999 = 10'h3cf == io_addr ? mem_975 : _GEN_1998; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2000 = 10'h3d0 == io_addr ? mem_976 : _GEN_1999; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2001 = 10'h3d1 == io_addr ? mem_977 : _GEN_2000; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2002 = 10'h3d2 == io_addr ? mem_978 : _GEN_2001; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2003 = 10'h3d3 == io_addr ? mem_979 : _GEN_2002; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2004 = 10'h3d4 == io_addr ? mem_980 : _GEN_2003; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2005 = 10'h3d5 == io_addr ? mem_981 : _GEN_2004; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2006 = 10'h3d6 == io_addr ? mem_982 : _GEN_2005; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2007 = 10'h3d7 == io_addr ? mem_983 : _GEN_2006; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2008 = 10'h3d8 == io_addr ? mem_984 : _GEN_2007; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2009 = 10'h3d9 == io_addr ? mem_985 : _GEN_2008; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2010 = 10'h3da == io_addr ? mem_986 : _GEN_2009; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2011 = 10'h3db == io_addr ? mem_987 : _GEN_2010; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2012 = 10'h3dc == io_addr ? mem_988 : _GEN_2011; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2013 = 10'h3dd == io_addr ? mem_989 : _GEN_2012; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2014 = 10'h3de == io_addr ? mem_990 : _GEN_2013; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2015 = 10'h3df == io_addr ? mem_991 : _GEN_2014; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2016 = 10'h3e0 == io_addr ? mem_992 : _GEN_2015; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2017 = 10'h3e1 == io_addr ? mem_993 : _GEN_2016; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2018 = 10'h3e2 == io_addr ? mem_994 : _GEN_2017; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2019 = 10'h3e3 == io_addr ? mem_995 : _GEN_2018; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2020 = 10'h3e4 == io_addr ? mem_996 : _GEN_2019; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2021 = 10'h3e5 == io_addr ? mem_997 : _GEN_2020; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2022 = 10'h3e6 == io_addr ? mem_998 : _GEN_2021; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2023 = 10'h3e7 == io_addr ? mem_999 : _GEN_2022; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2024 = 10'h3e8 == io_addr ? mem_1000 : _GEN_2023; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2025 = 10'h3e9 == io_addr ? mem_1001 : _GEN_2024; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2026 = 10'h3ea == io_addr ? mem_1002 : _GEN_2025; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2027 = 10'h3eb == io_addr ? mem_1003 : _GEN_2026; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2028 = 10'h3ec == io_addr ? mem_1004 : _GEN_2027; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2029 = 10'h3ed == io_addr ? mem_1005 : _GEN_2028; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2030 = 10'h3ee == io_addr ? mem_1006 : _GEN_2029; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2031 = 10'h3ef == io_addr ? mem_1007 : _GEN_2030; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2032 = 10'h3f0 == io_addr ? mem_1008 : _GEN_2031; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2033 = 10'h3f1 == io_addr ? mem_1009 : _GEN_2032; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2034 = 10'h3f2 == io_addr ? mem_1010 : _GEN_2033; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2035 = 10'h3f3 == io_addr ? mem_1011 : _GEN_2034; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2036 = 10'h3f4 == io_addr ? mem_1012 : _GEN_2035; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2037 = 10'h3f5 == io_addr ? mem_1013 : _GEN_2036; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2038 = 10'h3f6 == io_addr ? mem_1014 : _GEN_2037; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2039 = 10'h3f7 == io_addr ? mem_1015 : _GEN_2038; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2040 = 10'h3f8 == io_addr ? mem_1016 : _GEN_2039; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2041 = 10'h3f9 == io_addr ? mem_1017 : _GEN_2040; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2042 = 10'h3fa == io_addr ? mem_1018 : _GEN_2041; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2043 = 10'h3fb == io_addr ? mem_1019 : _GEN_2042; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2044 = 10'h3fc == io_addr ? mem_1020 : _GEN_2043; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2045 = 10'h3fd == io_addr ? mem_1021 : _GEN_2044; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2046 = 10'h3fe == io_addr ? mem_1022 : _GEN_2045; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_2047 = 10'h3ff == io_addr ? mem_1023 : _GEN_2046; // @[Ram.scala 20:{31,31}]
  wire [255:0] _GEN_3072 = io_write ? 256'h0 : _GEN_2047; // @[Ram.scala 17:14 19:20 20:31]
  assign io_dataOut = io_enable ? _GEN_3072 : 256'h0; // @[Ram.scala 17:14 18:19]
  always @(posedge clock) begin
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h0 == io_addr) begin // @[Ram.scala 19:35]
          mem_0 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1 == io_addr) begin // @[Ram.scala 19:35]
          mem_1 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2 == io_addr) begin // @[Ram.scala 19:35]
          mem_2 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3 == io_addr) begin // @[Ram.scala 19:35]
          mem_3 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h4 == io_addr) begin // @[Ram.scala 19:35]
          mem_4 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h5 == io_addr) begin // @[Ram.scala 19:35]
          mem_5 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h6 == io_addr) begin // @[Ram.scala 19:35]
          mem_6 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h7 == io_addr) begin // @[Ram.scala 19:35]
          mem_7 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h8 == io_addr) begin // @[Ram.scala 19:35]
          mem_8 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h9 == io_addr) begin // @[Ram.scala 19:35]
          mem_9 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'ha == io_addr) begin // @[Ram.scala 19:35]
          mem_10 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hb == io_addr) begin // @[Ram.scala 19:35]
          mem_11 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hc == io_addr) begin // @[Ram.scala 19:35]
          mem_12 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hd == io_addr) begin // @[Ram.scala 19:35]
          mem_13 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'he == io_addr) begin // @[Ram.scala 19:35]
          mem_14 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hf == io_addr) begin // @[Ram.scala 19:35]
          mem_15 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h10 == io_addr) begin // @[Ram.scala 19:35]
          mem_16 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h11 == io_addr) begin // @[Ram.scala 19:35]
          mem_17 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h12 == io_addr) begin // @[Ram.scala 19:35]
          mem_18 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h13 == io_addr) begin // @[Ram.scala 19:35]
          mem_19 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h14 == io_addr) begin // @[Ram.scala 19:35]
          mem_20 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h15 == io_addr) begin // @[Ram.scala 19:35]
          mem_21 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h16 == io_addr) begin // @[Ram.scala 19:35]
          mem_22 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h17 == io_addr) begin // @[Ram.scala 19:35]
          mem_23 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h18 == io_addr) begin // @[Ram.scala 19:35]
          mem_24 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h19 == io_addr) begin // @[Ram.scala 19:35]
          mem_25 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1a == io_addr) begin // @[Ram.scala 19:35]
          mem_26 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1b == io_addr) begin // @[Ram.scala 19:35]
          mem_27 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1c == io_addr) begin // @[Ram.scala 19:35]
          mem_28 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1d == io_addr) begin // @[Ram.scala 19:35]
          mem_29 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1e == io_addr) begin // @[Ram.scala 19:35]
          mem_30 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1f == io_addr) begin // @[Ram.scala 19:35]
          mem_31 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h20 == io_addr) begin // @[Ram.scala 19:35]
          mem_32 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h21 == io_addr) begin // @[Ram.scala 19:35]
          mem_33 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h22 == io_addr) begin // @[Ram.scala 19:35]
          mem_34 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h23 == io_addr) begin // @[Ram.scala 19:35]
          mem_35 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h24 == io_addr) begin // @[Ram.scala 19:35]
          mem_36 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h25 == io_addr) begin // @[Ram.scala 19:35]
          mem_37 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h26 == io_addr) begin // @[Ram.scala 19:35]
          mem_38 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h27 == io_addr) begin // @[Ram.scala 19:35]
          mem_39 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h28 == io_addr) begin // @[Ram.scala 19:35]
          mem_40 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h29 == io_addr) begin // @[Ram.scala 19:35]
          mem_41 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2a == io_addr) begin // @[Ram.scala 19:35]
          mem_42 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2b == io_addr) begin // @[Ram.scala 19:35]
          mem_43 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2c == io_addr) begin // @[Ram.scala 19:35]
          mem_44 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2d == io_addr) begin // @[Ram.scala 19:35]
          mem_45 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2e == io_addr) begin // @[Ram.scala 19:35]
          mem_46 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2f == io_addr) begin // @[Ram.scala 19:35]
          mem_47 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h30 == io_addr) begin // @[Ram.scala 19:35]
          mem_48 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h31 == io_addr) begin // @[Ram.scala 19:35]
          mem_49 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h32 == io_addr) begin // @[Ram.scala 19:35]
          mem_50 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h33 == io_addr) begin // @[Ram.scala 19:35]
          mem_51 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h34 == io_addr) begin // @[Ram.scala 19:35]
          mem_52 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h35 == io_addr) begin // @[Ram.scala 19:35]
          mem_53 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h36 == io_addr) begin // @[Ram.scala 19:35]
          mem_54 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h37 == io_addr) begin // @[Ram.scala 19:35]
          mem_55 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h38 == io_addr) begin // @[Ram.scala 19:35]
          mem_56 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h39 == io_addr) begin // @[Ram.scala 19:35]
          mem_57 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3a == io_addr) begin // @[Ram.scala 19:35]
          mem_58 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3b == io_addr) begin // @[Ram.scala 19:35]
          mem_59 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3c == io_addr) begin // @[Ram.scala 19:35]
          mem_60 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3d == io_addr) begin // @[Ram.scala 19:35]
          mem_61 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3e == io_addr) begin // @[Ram.scala 19:35]
          mem_62 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3f == io_addr) begin // @[Ram.scala 19:35]
          mem_63 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h40 == io_addr) begin // @[Ram.scala 19:35]
          mem_64 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h41 == io_addr) begin // @[Ram.scala 19:35]
          mem_65 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h42 == io_addr) begin // @[Ram.scala 19:35]
          mem_66 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h43 == io_addr) begin // @[Ram.scala 19:35]
          mem_67 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h44 == io_addr) begin // @[Ram.scala 19:35]
          mem_68 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h45 == io_addr) begin // @[Ram.scala 19:35]
          mem_69 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h46 == io_addr) begin // @[Ram.scala 19:35]
          mem_70 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h47 == io_addr) begin // @[Ram.scala 19:35]
          mem_71 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h48 == io_addr) begin // @[Ram.scala 19:35]
          mem_72 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h49 == io_addr) begin // @[Ram.scala 19:35]
          mem_73 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h4a == io_addr) begin // @[Ram.scala 19:35]
          mem_74 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h4b == io_addr) begin // @[Ram.scala 19:35]
          mem_75 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h4c == io_addr) begin // @[Ram.scala 19:35]
          mem_76 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h4d == io_addr) begin // @[Ram.scala 19:35]
          mem_77 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h4e == io_addr) begin // @[Ram.scala 19:35]
          mem_78 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h4f == io_addr) begin // @[Ram.scala 19:35]
          mem_79 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h50 == io_addr) begin // @[Ram.scala 19:35]
          mem_80 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h51 == io_addr) begin // @[Ram.scala 19:35]
          mem_81 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h52 == io_addr) begin // @[Ram.scala 19:35]
          mem_82 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h53 == io_addr) begin // @[Ram.scala 19:35]
          mem_83 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h54 == io_addr) begin // @[Ram.scala 19:35]
          mem_84 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h55 == io_addr) begin // @[Ram.scala 19:35]
          mem_85 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h56 == io_addr) begin // @[Ram.scala 19:35]
          mem_86 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h57 == io_addr) begin // @[Ram.scala 19:35]
          mem_87 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h58 == io_addr) begin // @[Ram.scala 19:35]
          mem_88 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h59 == io_addr) begin // @[Ram.scala 19:35]
          mem_89 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h5a == io_addr) begin // @[Ram.scala 19:35]
          mem_90 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h5b == io_addr) begin // @[Ram.scala 19:35]
          mem_91 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h5c == io_addr) begin // @[Ram.scala 19:35]
          mem_92 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h5d == io_addr) begin // @[Ram.scala 19:35]
          mem_93 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h5e == io_addr) begin // @[Ram.scala 19:35]
          mem_94 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h5f == io_addr) begin // @[Ram.scala 19:35]
          mem_95 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h60 == io_addr) begin // @[Ram.scala 19:35]
          mem_96 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h61 == io_addr) begin // @[Ram.scala 19:35]
          mem_97 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h62 == io_addr) begin // @[Ram.scala 19:35]
          mem_98 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h63 == io_addr) begin // @[Ram.scala 19:35]
          mem_99 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h64 == io_addr) begin // @[Ram.scala 19:35]
          mem_100 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h65 == io_addr) begin // @[Ram.scala 19:35]
          mem_101 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h66 == io_addr) begin // @[Ram.scala 19:35]
          mem_102 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h67 == io_addr) begin // @[Ram.scala 19:35]
          mem_103 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h68 == io_addr) begin // @[Ram.scala 19:35]
          mem_104 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h69 == io_addr) begin // @[Ram.scala 19:35]
          mem_105 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h6a == io_addr) begin // @[Ram.scala 19:35]
          mem_106 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h6b == io_addr) begin // @[Ram.scala 19:35]
          mem_107 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h6c == io_addr) begin // @[Ram.scala 19:35]
          mem_108 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h6d == io_addr) begin // @[Ram.scala 19:35]
          mem_109 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h6e == io_addr) begin // @[Ram.scala 19:35]
          mem_110 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h6f == io_addr) begin // @[Ram.scala 19:35]
          mem_111 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h70 == io_addr) begin // @[Ram.scala 19:35]
          mem_112 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h71 == io_addr) begin // @[Ram.scala 19:35]
          mem_113 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h72 == io_addr) begin // @[Ram.scala 19:35]
          mem_114 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h73 == io_addr) begin // @[Ram.scala 19:35]
          mem_115 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h74 == io_addr) begin // @[Ram.scala 19:35]
          mem_116 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h75 == io_addr) begin // @[Ram.scala 19:35]
          mem_117 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h76 == io_addr) begin // @[Ram.scala 19:35]
          mem_118 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h77 == io_addr) begin // @[Ram.scala 19:35]
          mem_119 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h78 == io_addr) begin // @[Ram.scala 19:35]
          mem_120 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h79 == io_addr) begin // @[Ram.scala 19:35]
          mem_121 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h7a == io_addr) begin // @[Ram.scala 19:35]
          mem_122 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h7b == io_addr) begin // @[Ram.scala 19:35]
          mem_123 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h7c == io_addr) begin // @[Ram.scala 19:35]
          mem_124 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h7d == io_addr) begin // @[Ram.scala 19:35]
          mem_125 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h7e == io_addr) begin // @[Ram.scala 19:35]
          mem_126 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h7f == io_addr) begin // @[Ram.scala 19:35]
          mem_127 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h80 == io_addr) begin // @[Ram.scala 19:35]
          mem_128 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h81 == io_addr) begin // @[Ram.scala 19:35]
          mem_129 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h82 == io_addr) begin // @[Ram.scala 19:35]
          mem_130 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h83 == io_addr) begin // @[Ram.scala 19:35]
          mem_131 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h84 == io_addr) begin // @[Ram.scala 19:35]
          mem_132 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h85 == io_addr) begin // @[Ram.scala 19:35]
          mem_133 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h86 == io_addr) begin // @[Ram.scala 19:35]
          mem_134 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h87 == io_addr) begin // @[Ram.scala 19:35]
          mem_135 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h88 == io_addr) begin // @[Ram.scala 19:35]
          mem_136 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h89 == io_addr) begin // @[Ram.scala 19:35]
          mem_137 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h8a == io_addr) begin // @[Ram.scala 19:35]
          mem_138 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h8b == io_addr) begin // @[Ram.scala 19:35]
          mem_139 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h8c == io_addr) begin // @[Ram.scala 19:35]
          mem_140 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h8d == io_addr) begin // @[Ram.scala 19:35]
          mem_141 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h8e == io_addr) begin // @[Ram.scala 19:35]
          mem_142 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h8f == io_addr) begin // @[Ram.scala 19:35]
          mem_143 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h90 == io_addr) begin // @[Ram.scala 19:35]
          mem_144 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h91 == io_addr) begin // @[Ram.scala 19:35]
          mem_145 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h92 == io_addr) begin // @[Ram.scala 19:35]
          mem_146 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h93 == io_addr) begin // @[Ram.scala 19:35]
          mem_147 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h94 == io_addr) begin // @[Ram.scala 19:35]
          mem_148 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h95 == io_addr) begin // @[Ram.scala 19:35]
          mem_149 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h96 == io_addr) begin // @[Ram.scala 19:35]
          mem_150 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h97 == io_addr) begin // @[Ram.scala 19:35]
          mem_151 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h98 == io_addr) begin // @[Ram.scala 19:35]
          mem_152 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h99 == io_addr) begin // @[Ram.scala 19:35]
          mem_153 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h9a == io_addr) begin // @[Ram.scala 19:35]
          mem_154 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h9b == io_addr) begin // @[Ram.scala 19:35]
          mem_155 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h9c == io_addr) begin // @[Ram.scala 19:35]
          mem_156 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h9d == io_addr) begin // @[Ram.scala 19:35]
          mem_157 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h9e == io_addr) begin // @[Ram.scala 19:35]
          mem_158 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h9f == io_addr) begin // @[Ram.scala 19:35]
          mem_159 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'ha0 == io_addr) begin // @[Ram.scala 19:35]
          mem_160 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'ha1 == io_addr) begin // @[Ram.scala 19:35]
          mem_161 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'ha2 == io_addr) begin // @[Ram.scala 19:35]
          mem_162 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'ha3 == io_addr) begin // @[Ram.scala 19:35]
          mem_163 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'ha4 == io_addr) begin // @[Ram.scala 19:35]
          mem_164 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'ha5 == io_addr) begin // @[Ram.scala 19:35]
          mem_165 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'ha6 == io_addr) begin // @[Ram.scala 19:35]
          mem_166 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'ha7 == io_addr) begin // @[Ram.scala 19:35]
          mem_167 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'ha8 == io_addr) begin // @[Ram.scala 19:35]
          mem_168 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'ha9 == io_addr) begin // @[Ram.scala 19:35]
          mem_169 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'haa == io_addr) begin // @[Ram.scala 19:35]
          mem_170 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hab == io_addr) begin // @[Ram.scala 19:35]
          mem_171 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hac == io_addr) begin // @[Ram.scala 19:35]
          mem_172 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'had == io_addr) begin // @[Ram.scala 19:35]
          mem_173 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hae == io_addr) begin // @[Ram.scala 19:35]
          mem_174 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'haf == io_addr) begin // @[Ram.scala 19:35]
          mem_175 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hb0 == io_addr) begin // @[Ram.scala 19:35]
          mem_176 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hb1 == io_addr) begin // @[Ram.scala 19:35]
          mem_177 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hb2 == io_addr) begin // @[Ram.scala 19:35]
          mem_178 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hb3 == io_addr) begin // @[Ram.scala 19:35]
          mem_179 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hb4 == io_addr) begin // @[Ram.scala 19:35]
          mem_180 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hb5 == io_addr) begin // @[Ram.scala 19:35]
          mem_181 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hb6 == io_addr) begin // @[Ram.scala 19:35]
          mem_182 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hb7 == io_addr) begin // @[Ram.scala 19:35]
          mem_183 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hb8 == io_addr) begin // @[Ram.scala 19:35]
          mem_184 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hb9 == io_addr) begin // @[Ram.scala 19:35]
          mem_185 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hba == io_addr) begin // @[Ram.scala 19:35]
          mem_186 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hbb == io_addr) begin // @[Ram.scala 19:35]
          mem_187 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hbc == io_addr) begin // @[Ram.scala 19:35]
          mem_188 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hbd == io_addr) begin // @[Ram.scala 19:35]
          mem_189 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hbe == io_addr) begin // @[Ram.scala 19:35]
          mem_190 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hbf == io_addr) begin // @[Ram.scala 19:35]
          mem_191 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hc0 == io_addr) begin // @[Ram.scala 19:35]
          mem_192 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hc1 == io_addr) begin // @[Ram.scala 19:35]
          mem_193 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hc2 == io_addr) begin // @[Ram.scala 19:35]
          mem_194 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hc3 == io_addr) begin // @[Ram.scala 19:35]
          mem_195 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hc4 == io_addr) begin // @[Ram.scala 19:35]
          mem_196 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hc5 == io_addr) begin // @[Ram.scala 19:35]
          mem_197 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hc6 == io_addr) begin // @[Ram.scala 19:35]
          mem_198 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hc7 == io_addr) begin // @[Ram.scala 19:35]
          mem_199 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hc8 == io_addr) begin // @[Ram.scala 19:35]
          mem_200 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hc9 == io_addr) begin // @[Ram.scala 19:35]
          mem_201 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hca == io_addr) begin // @[Ram.scala 19:35]
          mem_202 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hcb == io_addr) begin // @[Ram.scala 19:35]
          mem_203 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hcc == io_addr) begin // @[Ram.scala 19:35]
          mem_204 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hcd == io_addr) begin // @[Ram.scala 19:35]
          mem_205 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hce == io_addr) begin // @[Ram.scala 19:35]
          mem_206 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hcf == io_addr) begin // @[Ram.scala 19:35]
          mem_207 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hd0 == io_addr) begin // @[Ram.scala 19:35]
          mem_208 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hd1 == io_addr) begin // @[Ram.scala 19:35]
          mem_209 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hd2 == io_addr) begin // @[Ram.scala 19:35]
          mem_210 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hd3 == io_addr) begin // @[Ram.scala 19:35]
          mem_211 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hd4 == io_addr) begin // @[Ram.scala 19:35]
          mem_212 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hd5 == io_addr) begin // @[Ram.scala 19:35]
          mem_213 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hd6 == io_addr) begin // @[Ram.scala 19:35]
          mem_214 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hd7 == io_addr) begin // @[Ram.scala 19:35]
          mem_215 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hd8 == io_addr) begin // @[Ram.scala 19:35]
          mem_216 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hd9 == io_addr) begin // @[Ram.scala 19:35]
          mem_217 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hda == io_addr) begin // @[Ram.scala 19:35]
          mem_218 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hdb == io_addr) begin // @[Ram.scala 19:35]
          mem_219 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hdc == io_addr) begin // @[Ram.scala 19:35]
          mem_220 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hdd == io_addr) begin // @[Ram.scala 19:35]
          mem_221 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hde == io_addr) begin // @[Ram.scala 19:35]
          mem_222 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hdf == io_addr) begin // @[Ram.scala 19:35]
          mem_223 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'he0 == io_addr) begin // @[Ram.scala 19:35]
          mem_224 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'he1 == io_addr) begin // @[Ram.scala 19:35]
          mem_225 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'he2 == io_addr) begin // @[Ram.scala 19:35]
          mem_226 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'he3 == io_addr) begin // @[Ram.scala 19:35]
          mem_227 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'he4 == io_addr) begin // @[Ram.scala 19:35]
          mem_228 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'he5 == io_addr) begin // @[Ram.scala 19:35]
          mem_229 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'he6 == io_addr) begin // @[Ram.scala 19:35]
          mem_230 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'he7 == io_addr) begin // @[Ram.scala 19:35]
          mem_231 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'he8 == io_addr) begin // @[Ram.scala 19:35]
          mem_232 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'he9 == io_addr) begin // @[Ram.scala 19:35]
          mem_233 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hea == io_addr) begin // @[Ram.scala 19:35]
          mem_234 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'heb == io_addr) begin // @[Ram.scala 19:35]
          mem_235 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hec == io_addr) begin // @[Ram.scala 19:35]
          mem_236 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hed == io_addr) begin // @[Ram.scala 19:35]
          mem_237 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hee == io_addr) begin // @[Ram.scala 19:35]
          mem_238 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hef == io_addr) begin // @[Ram.scala 19:35]
          mem_239 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hf0 == io_addr) begin // @[Ram.scala 19:35]
          mem_240 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hf1 == io_addr) begin // @[Ram.scala 19:35]
          mem_241 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hf2 == io_addr) begin // @[Ram.scala 19:35]
          mem_242 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hf3 == io_addr) begin // @[Ram.scala 19:35]
          mem_243 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hf4 == io_addr) begin // @[Ram.scala 19:35]
          mem_244 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hf5 == io_addr) begin // @[Ram.scala 19:35]
          mem_245 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hf6 == io_addr) begin // @[Ram.scala 19:35]
          mem_246 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hf7 == io_addr) begin // @[Ram.scala 19:35]
          mem_247 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hf8 == io_addr) begin // @[Ram.scala 19:35]
          mem_248 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hf9 == io_addr) begin // @[Ram.scala 19:35]
          mem_249 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hfa == io_addr) begin // @[Ram.scala 19:35]
          mem_250 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hfb == io_addr) begin // @[Ram.scala 19:35]
          mem_251 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hfc == io_addr) begin // @[Ram.scala 19:35]
          mem_252 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hfd == io_addr) begin // @[Ram.scala 19:35]
          mem_253 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hfe == io_addr) begin // @[Ram.scala 19:35]
          mem_254 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'hff == io_addr) begin // @[Ram.scala 19:35]
          mem_255 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h100 == io_addr) begin // @[Ram.scala 19:35]
          mem_256 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h101 == io_addr) begin // @[Ram.scala 19:35]
          mem_257 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h102 == io_addr) begin // @[Ram.scala 19:35]
          mem_258 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h103 == io_addr) begin // @[Ram.scala 19:35]
          mem_259 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h104 == io_addr) begin // @[Ram.scala 19:35]
          mem_260 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h105 == io_addr) begin // @[Ram.scala 19:35]
          mem_261 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h106 == io_addr) begin // @[Ram.scala 19:35]
          mem_262 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h107 == io_addr) begin // @[Ram.scala 19:35]
          mem_263 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h108 == io_addr) begin // @[Ram.scala 19:35]
          mem_264 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h109 == io_addr) begin // @[Ram.scala 19:35]
          mem_265 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h10a == io_addr) begin // @[Ram.scala 19:35]
          mem_266 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h10b == io_addr) begin // @[Ram.scala 19:35]
          mem_267 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h10c == io_addr) begin // @[Ram.scala 19:35]
          mem_268 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h10d == io_addr) begin // @[Ram.scala 19:35]
          mem_269 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h10e == io_addr) begin // @[Ram.scala 19:35]
          mem_270 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h10f == io_addr) begin // @[Ram.scala 19:35]
          mem_271 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h110 == io_addr) begin // @[Ram.scala 19:35]
          mem_272 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h111 == io_addr) begin // @[Ram.scala 19:35]
          mem_273 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h112 == io_addr) begin // @[Ram.scala 19:35]
          mem_274 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h113 == io_addr) begin // @[Ram.scala 19:35]
          mem_275 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h114 == io_addr) begin // @[Ram.scala 19:35]
          mem_276 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h115 == io_addr) begin // @[Ram.scala 19:35]
          mem_277 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h116 == io_addr) begin // @[Ram.scala 19:35]
          mem_278 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h117 == io_addr) begin // @[Ram.scala 19:35]
          mem_279 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h118 == io_addr) begin // @[Ram.scala 19:35]
          mem_280 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h119 == io_addr) begin // @[Ram.scala 19:35]
          mem_281 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h11a == io_addr) begin // @[Ram.scala 19:35]
          mem_282 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h11b == io_addr) begin // @[Ram.scala 19:35]
          mem_283 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h11c == io_addr) begin // @[Ram.scala 19:35]
          mem_284 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h11d == io_addr) begin // @[Ram.scala 19:35]
          mem_285 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h11e == io_addr) begin // @[Ram.scala 19:35]
          mem_286 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h11f == io_addr) begin // @[Ram.scala 19:35]
          mem_287 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h120 == io_addr) begin // @[Ram.scala 19:35]
          mem_288 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h121 == io_addr) begin // @[Ram.scala 19:35]
          mem_289 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h122 == io_addr) begin // @[Ram.scala 19:35]
          mem_290 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h123 == io_addr) begin // @[Ram.scala 19:35]
          mem_291 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h124 == io_addr) begin // @[Ram.scala 19:35]
          mem_292 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h125 == io_addr) begin // @[Ram.scala 19:35]
          mem_293 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h126 == io_addr) begin // @[Ram.scala 19:35]
          mem_294 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h127 == io_addr) begin // @[Ram.scala 19:35]
          mem_295 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h128 == io_addr) begin // @[Ram.scala 19:35]
          mem_296 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h129 == io_addr) begin // @[Ram.scala 19:35]
          mem_297 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h12a == io_addr) begin // @[Ram.scala 19:35]
          mem_298 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h12b == io_addr) begin // @[Ram.scala 19:35]
          mem_299 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h12c == io_addr) begin // @[Ram.scala 19:35]
          mem_300 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h12d == io_addr) begin // @[Ram.scala 19:35]
          mem_301 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h12e == io_addr) begin // @[Ram.scala 19:35]
          mem_302 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h12f == io_addr) begin // @[Ram.scala 19:35]
          mem_303 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h130 == io_addr) begin // @[Ram.scala 19:35]
          mem_304 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h131 == io_addr) begin // @[Ram.scala 19:35]
          mem_305 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h132 == io_addr) begin // @[Ram.scala 19:35]
          mem_306 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h133 == io_addr) begin // @[Ram.scala 19:35]
          mem_307 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h134 == io_addr) begin // @[Ram.scala 19:35]
          mem_308 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h135 == io_addr) begin // @[Ram.scala 19:35]
          mem_309 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h136 == io_addr) begin // @[Ram.scala 19:35]
          mem_310 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h137 == io_addr) begin // @[Ram.scala 19:35]
          mem_311 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h138 == io_addr) begin // @[Ram.scala 19:35]
          mem_312 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h139 == io_addr) begin // @[Ram.scala 19:35]
          mem_313 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h13a == io_addr) begin // @[Ram.scala 19:35]
          mem_314 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h13b == io_addr) begin // @[Ram.scala 19:35]
          mem_315 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h13c == io_addr) begin // @[Ram.scala 19:35]
          mem_316 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h13d == io_addr) begin // @[Ram.scala 19:35]
          mem_317 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h13e == io_addr) begin // @[Ram.scala 19:35]
          mem_318 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h13f == io_addr) begin // @[Ram.scala 19:35]
          mem_319 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h140 == io_addr) begin // @[Ram.scala 19:35]
          mem_320 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h141 == io_addr) begin // @[Ram.scala 19:35]
          mem_321 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h142 == io_addr) begin // @[Ram.scala 19:35]
          mem_322 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h143 == io_addr) begin // @[Ram.scala 19:35]
          mem_323 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h144 == io_addr) begin // @[Ram.scala 19:35]
          mem_324 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h145 == io_addr) begin // @[Ram.scala 19:35]
          mem_325 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h146 == io_addr) begin // @[Ram.scala 19:35]
          mem_326 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h147 == io_addr) begin // @[Ram.scala 19:35]
          mem_327 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h148 == io_addr) begin // @[Ram.scala 19:35]
          mem_328 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h149 == io_addr) begin // @[Ram.scala 19:35]
          mem_329 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h14a == io_addr) begin // @[Ram.scala 19:35]
          mem_330 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h14b == io_addr) begin // @[Ram.scala 19:35]
          mem_331 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h14c == io_addr) begin // @[Ram.scala 19:35]
          mem_332 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h14d == io_addr) begin // @[Ram.scala 19:35]
          mem_333 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h14e == io_addr) begin // @[Ram.scala 19:35]
          mem_334 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h14f == io_addr) begin // @[Ram.scala 19:35]
          mem_335 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h150 == io_addr) begin // @[Ram.scala 19:35]
          mem_336 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h151 == io_addr) begin // @[Ram.scala 19:35]
          mem_337 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h152 == io_addr) begin // @[Ram.scala 19:35]
          mem_338 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h153 == io_addr) begin // @[Ram.scala 19:35]
          mem_339 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h154 == io_addr) begin // @[Ram.scala 19:35]
          mem_340 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h155 == io_addr) begin // @[Ram.scala 19:35]
          mem_341 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h156 == io_addr) begin // @[Ram.scala 19:35]
          mem_342 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h157 == io_addr) begin // @[Ram.scala 19:35]
          mem_343 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h158 == io_addr) begin // @[Ram.scala 19:35]
          mem_344 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h159 == io_addr) begin // @[Ram.scala 19:35]
          mem_345 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h15a == io_addr) begin // @[Ram.scala 19:35]
          mem_346 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h15b == io_addr) begin // @[Ram.scala 19:35]
          mem_347 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h15c == io_addr) begin // @[Ram.scala 19:35]
          mem_348 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h15d == io_addr) begin // @[Ram.scala 19:35]
          mem_349 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h15e == io_addr) begin // @[Ram.scala 19:35]
          mem_350 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h15f == io_addr) begin // @[Ram.scala 19:35]
          mem_351 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h160 == io_addr) begin // @[Ram.scala 19:35]
          mem_352 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h161 == io_addr) begin // @[Ram.scala 19:35]
          mem_353 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h162 == io_addr) begin // @[Ram.scala 19:35]
          mem_354 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h163 == io_addr) begin // @[Ram.scala 19:35]
          mem_355 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h164 == io_addr) begin // @[Ram.scala 19:35]
          mem_356 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h165 == io_addr) begin // @[Ram.scala 19:35]
          mem_357 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h166 == io_addr) begin // @[Ram.scala 19:35]
          mem_358 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h167 == io_addr) begin // @[Ram.scala 19:35]
          mem_359 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h168 == io_addr) begin // @[Ram.scala 19:35]
          mem_360 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h169 == io_addr) begin // @[Ram.scala 19:35]
          mem_361 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h16a == io_addr) begin // @[Ram.scala 19:35]
          mem_362 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h16b == io_addr) begin // @[Ram.scala 19:35]
          mem_363 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h16c == io_addr) begin // @[Ram.scala 19:35]
          mem_364 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h16d == io_addr) begin // @[Ram.scala 19:35]
          mem_365 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h16e == io_addr) begin // @[Ram.scala 19:35]
          mem_366 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h16f == io_addr) begin // @[Ram.scala 19:35]
          mem_367 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h170 == io_addr) begin // @[Ram.scala 19:35]
          mem_368 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h171 == io_addr) begin // @[Ram.scala 19:35]
          mem_369 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h172 == io_addr) begin // @[Ram.scala 19:35]
          mem_370 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h173 == io_addr) begin // @[Ram.scala 19:35]
          mem_371 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h174 == io_addr) begin // @[Ram.scala 19:35]
          mem_372 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h175 == io_addr) begin // @[Ram.scala 19:35]
          mem_373 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h176 == io_addr) begin // @[Ram.scala 19:35]
          mem_374 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h177 == io_addr) begin // @[Ram.scala 19:35]
          mem_375 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h178 == io_addr) begin // @[Ram.scala 19:35]
          mem_376 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h179 == io_addr) begin // @[Ram.scala 19:35]
          mem_377 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h17a == io_addr) begin // @[Ram.scala 19:35]
          mem_378 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h17b == io_addr) begin // @[Ram.scala 19:35]
          mem_379 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h17c == io_addr) begin // @[Ram.scala 19:35]
          mem_380 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h17d == io_addr) begin // @[Ram.scala 19:35]
          mem_381 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h17e == io_addr) begin // @[Ram.scala 19:35]
          mem_382 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h17f == io_addr) begin // @[Ram.scala 19:35]
          mem_383 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h180 == io_addr) begin // @[Ram.scala 19:35]
          mem_384 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h181 == io_addr) begin // @[Ram.scala 19:35]
          mem_385 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h182 == io_addr) begin // @[Ram.scala 19:35]
          mem_386 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h183 == io_addr) begin // @[Ram.scala 19:35]
          mem_387 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h184 == io_addr) begin // @[Ram.scala 19:35]
          mem_388 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h185 == io_addr) begin // @[Ram.scala 19:35]
          mem_389 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h186 == io_addr) begin // @[Ram.scala 19:35]
          mem_390 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h187 == io_addr) begin // @[Ram.scala 19:35]
          mem_391 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h188 == io_addr) begin // @[Ram.scala 19:35]
          mem_392 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h189 == io_addr) begin // @[Ram.scala 19:35]
          mem_393 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h18a == io_addr) begin // @[Ram.scala 19:35]
          mem_394 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h18b == io_addr) begin // @[Ram.scala 19:35]
          mem_395 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h18c == io_addr) begin // @[Ram.scala 19:35]
          mem_396 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h18d == io_addr) begin // @[Ram.scala 19:35]
          mem_397 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h18e == io_addr) begin // @[Ram.scala 19:35]
          mem_398 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h18f == io_addr) begin // @[Ram.scala 19:35]
          mem_399 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h190 == io_addr) begin // @[Ram.scala 19:35]
          mem_400 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h191 == io_addr) begin // @[Ram.scala 19:35]
          mem_401 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h192 == io_addr) begin // @[Ram.scala 19:35]
          mem_402 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h193 == io_addr) begin // @[Ram.scala 19:35]
          mem_403 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h194 == io_addr) begin // @[Ram.scala 19:35]
          mem_404 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h195 == io_addr) begin // @[Ram.scala 19:35]
          mem_405 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h196 == io_addr) begin // @[Ram.scala 19:35]
          mem_406 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h197 == io_addr) begin // @[Ram.scala 19:35]
          mem_407 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h198 == io_addr) begin // @[Ram.scala 19:35]
          mem_408 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h199 == io_addr) begin // @[Ram.scala 19:35]
          mem_409 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h19a == io_addr) begin // @[Ram.scala 19:35]
          mem_410 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h19b == io_addr) begin // @[Ram.scala 19:35]
          mem_411 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h19c == io_addr) begin // @[Ram.scala 19:35]
          mem_412 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h19d == io_addr) begin // @[Ram.scala 19:35]
          mem_413 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h19e == io_addr) begin // @[Ram.scala 19:35]
          mem_414 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h19f == io_addr) begin // @[Ram.scala 19:35]
          mem_415 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1a0 == io_addr) begin // @[Ram.scala 19:35]
          mem_416 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1a1 == io_addr) begin // @[Ram.scala 19:35]
          mem_417 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1a2 == io_addr) begin // @[Ram.scala 19:35]
          mem_418 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1a3 == io_addr) begin // @[Ram.scala 19:35]
          mem_419 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1a4 == io_addr) begin // @[Ram.scala 19:35]
          mem_420 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1a5 == io_addr) begin // @[Ram.scala 19:35]
          mem_421 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1a6 == io_addr) begin // @[Ram.scala 19:35]
          mem_422 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1a7 == io_addr) begin // @[Ram.scala 19:35]
          mem_423 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1a8 == io_addr) begin // @[Ram.scala 19:35]
          mem_424 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1a9 == io_addr) begin // @[Ram.scala 19:35]
          mem_425 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1aa == io_addr) begin // @[Ram.scala 19:35]
          mem_426 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ab == io_addr) begin // @[Ram.scala 19:35]
          mem_427 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ac == io_addr) begin // @[Ram.scala 19:35]
          mem_428 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ad == io_addr) begin // @[Ram.scala 19:35]
          mem_429 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ae == io_addr) begin // @[Ram.scala 19:35]
          mem_430 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1af == io_addr) begin // @[Ram.scala 19:35]
          mem_431 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1b0 == io_addr) begin // @[Ram.scala 19:35]
          mem_432 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1b1 == io_addr) begin // @[Ram.scala 19:35]
          mem_433 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1b2 == io_addr) begin // @[Ram.scala 19:35]
          mem_434 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1b3 == io_addr) begin // @[Ram.scala 19:35]
          mem_435 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1b4 == io_addr) begin // @[Ram.scala 19:35]
          mem_436 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1b5 == io_addr) begin // @[Ram.scala 19:35]
          mem_437 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1b6 == io_addr) begin // @[Ram.scala 19:35]
          mem_438 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1b7 == io_addr) begin // @[Ram.scala 19:35]
          mem_439 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1b8 == io_addr) begin // @[Ram.scala 19:35]
          mem_440 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1b9 == io_addr) begin // @[Ram.scala 19:35]
          mem_441 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ba == io_addr) begin // @[Ram.scala 19:35]
          mem_442 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1bb == io_addr) begin // @[Ram.scala 19:35]
          mem_443 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1bc == io_addr) begin // @[Ram.scala 19:35]
          mem_444 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1bd == io_addr) begin // @[Ram.scala 19:35]
          mem_445 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1be == io_addr) begin // @[Ram.scala 19:35]
          mem_446 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1bf == io_addr) begin // @[Ram.scala 19:35]
          mem_447 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1c0 == io_addr) begin // @[Ram.scala 19:35]
          mem_448 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1c1 == io_addr) begin // @[Ram.scala 19:35]
          mem_449 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1c2 == io_addr) begin // @[Ram.scala 19:35]
          mem_450 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1c3 == io_addr) begin // @[Ram.scala 19:35]
          mem_451 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1c4 == io_addr) begin // @[Ram.scala 19:35]
          mem_452 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1c5 == io_addr) begin // @[Ram.scala 19:35]
          mem_453 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1c6 == io_addr) begin // @[Ram.scala 19:35]
          mem_454 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1c7 == io_addr) begin // @[Ram.scala 19:35]
          mem_455 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1c8 == io_addr) begin // @[Ram.scala 19:35]
          mem_456 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1c9 == io_addr) begin // @[Ram.scala 19:35]
          mem_457 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ca == io_addr) begin // @[Ram.scala 19:35]
          mem_458 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1cb == io_addr) begin // @[Ram.scala 19:35]
          mem_459 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1cc == io_addr) begin // @[Ram.scala 19:35]
          mem_460 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1cd == io_addr) begin // @[Ram.scala 19:35]
          mem_461 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ce == io_addr) begin // @[Ram.scala 19:35]
          mem_462 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1cf == io_addr) begin // @[Ram.scala 19:35]
          mem_463 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1d0 == io_addr) begin // @[Ram.scala 19:35]
          mem_464 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1d1 == io_addr) begin // @[Ram.scala 19:35]
          mem_465 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1d2 == io_addr) begin // @[Ram.scala 19:35]
          mem_466 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1d3 == io_addr) begin // @[Ram.scala 19:35]
          mem_467 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1d4 == io_addr) begin // @[Ram.scala 19:35]
          mem_468 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1d5 == io_addr) begin // @[Ram.scala 19:35]
          mem_469 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1d6 == io_addr) begin // @[Ram.scala 19:35]
          mem_470 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1d7 == io_addr) begin // @[Ram.scala 19:35]
          mem_471 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1d8 == io_addr) begin // @[Ram.scala 19:35]
          mem_472 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1d9 == io_addr) begin // @[Ram.scala 19:35]
          mem_473 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1da == io_addr) begin // @[Ram.scala 19:35]
          mem_474 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1db == io_addr) begin // @[Ram.scala 19:35]
          mem_475 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1dc == io_addr) begin // @[Ram.scala 19:35]
          mem_476 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1dd == io_addr) begin // @[Ram.scala 19:35]
          mem_477 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1de == io_addr) begin // @[Ram.scala 19:35]
          mem_478 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1df == io_addr) begin // @[Ram.scala 19:35]
          mem_479 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1e0 == io_addr) begin // @[Ram.scala 19:35]
          mem_480 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1e1 == io_addr) begin // @[Ram.scala 19:35]
          mem_481 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1e2 == io_addr) begin // @[Ram.scala 19:35]
          mem_482 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1e3 == io_addr) begin // @[Ram.scala 19:35]
          mem_483 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1e4 == io_addr) begin // @[Ram.scala 19:35]
          mem_484 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1e5 == io_addr) begin // @[Ram.scala 19:35]
          mem_485 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1e6 == io_addr) begin // @[Ram.scala 19:35]
          mem_486 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1e7 == io_addr) begin // @[Ram.scala 19:35]
          mem_487 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1e8 == io_addr) begin // @[Ram.scala 19:35]
          mem_488 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1e9 == io_addr) begin // @[Ram.scala 19:35]
          mem_489 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ea == io_addr) begin // @[Ram.scala 19:35]
          mem_490 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1eb == io_addr) begin // @[Ram.scala 19:35]
          mem_491 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ec == io_addr) begin // @[Ram.scala 19:35]
          mem_492 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ed == io_addr) begin // @[Ram.scala 19:35]
          mem_493 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ee == io_addr) begin // @[Ram.scala 19:35]
          mem_494 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ef == io_addr) begin // @[Ram.scala 19:35]
          mem_495 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1f0 == io_addr) begin // @[Ram.scala 19:35]
          mem_496 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1f1 == io_addr) begin // @[Ram.scala 19:35]
          mem_497 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1f2 == io_addr) begin // @[Ram.scala 19:35]
          mem_498 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1f3 == io_addr) begin // @[Ram.scala 19:35]
          mem_499 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1f4 == io_addr) begin // @[Ram.scala 19:35]
          mem_500 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1f5 == io_addr) begin // @[Ram.scala 19:35]
          mem_501 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1f6 == io_addr) begin // @[Ram.scala 19:35]
          mem_502 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1f7 == io_addr) begin // @[Ram.scala 19:35]
          mem_503 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1f8 == io_addr) begin // @[Ram.scala 19:35]
          mem_504 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1f9 == io_addr) begin // @[Ram.scala 19:35]
          mem_505 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1fa == io_addr) begin // @[Ram.scala 19:35]
          mem_506 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1fb == io_addr) begin // @[Ram.scala 19:35]
          mem_507 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1fc == io_addr) begin // @[Ram.scala 19:35]
          mem_508 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1fd == io_addr) begin // @[Ram.scala 19:35]
          mem_509 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1fe == io_addr) begin // @[Ram.scala 19:35]
          mem_510 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h1ff == io_addr) begin // @[Ram.scala 19:35]
          mem_511 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h200 == io_addr) begin // @[Ram.scala 19:35]
          mem_512 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h201 == io_addr) begin // @[Ram.scala 19:35]
          mem_513 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h202 == io_addr) begin // @[Ram.scala 19:35]
          mem_514 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h203 == io_addr) begin // @[Ram.scala 19:35]
          mem_515 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h204 == io_addr) begin // @[Ram.scala 19:35]
          mem_516 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h205 == io_addr) begin // @[Ram.scala 19:35]
          mem_517 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h206 == io_addr) begin // @[Ram.scala 19:35]
          mem_518 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h207 == io_addr) begin // @[Ram.scala 19:35]
          mem_519 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h208 == io_addr) begin // @[Ram.scala 19:35]
          mem_520 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h209 == io_addr) begin // @[Ram.scala 19:35]
          mem_521 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h20a == io_addr) begin // @[Ram.scala 19:35]
          mem_522 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h20b == io_addr) begin // @[Ram.scala 19:35]
          mem_523 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h20c == io_addr) begin // @[Ram.scala 19:35]
          mem_524 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h20d == io_addr) begin // @[Ram.scala 19:35]
          mem_525 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h20e == io_addr) begin // @[Ram.scala 19:35]
          mem_526 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h20f == io_addr) begin // @[Ram.scala 19:35]
          mem_527 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h210 == io_addr) begin // @[Ram.scala 19:35]
          mem_528 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h211 == io_addr) begin // @[Ram.scala 19:35]
          mem_529 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h212 == io_addr) begin // @[Ram.scala 19:35]
          mem_530 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h213 == io_addr) begin // @[Ram.scala 19:35]
          mem_531 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h214 == io_addr) begin // @[Ram.scala 19:35]
          mem_532 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h215 == io_addr) begin // @[Ram.scala 19:35]
          mem_533 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h216 == io_addr) begin // @[Ram.scala 19:35]
          mem_534 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h217 == io_addr) begin // @[Ram.scala 19:35]
          mem_535 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h218 == io_addr) begin // @[Ram.scala 19:35]
          mem_536 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h219 == io_addr) begin // @[Ram.scala 19:35]
          mem_537 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h21a == io_addr) begin // @[Ram.scala 19:35]
          mem_538 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h21b == io_addr) begin // @[Ram.scala 19:35]
          mem_539 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h21c == io_addr) begin // @[Ram.scala 19:35]
          mem_540 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h21d == io_addr) begin // @[Ram.scala 19:35]
          mem_541 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h21e == io_addr) begin // @[Ram.scala 19:35]
          mem_542 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h21f == io_addr) begin // @[Ram.scala 19:35]
          mem_543 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h220 == io_addr) begin // @[Ram.scala 19:35]
          mem_544 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h221 == io_addr) begin // @[Ram.scala 19:35]
          mem_545 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h222 == io_addr) begin // @[Ram.scala 19:35]
          mem_546 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h223 == io_addr) begin // @[Ram.scala 19:35]
          mem_547 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h224 == io_addr) begin // @[Ram.scala 19:35]
          mem_548 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h225 == io_addr) begin // @[Ram.scala 19:35]
          mem_549 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h226 == io_addr) begin // @[Ram.scala 19:35]
          mem_550 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h227 == io_addr) begin // @[Ram.scala 19:35]
          mem_551 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h228 == io_addr) begin // @[Ram.scala 19:35]
          mem_552 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h229 == io_addr) begin // @[Ram.scala 19:35]
          mem_553 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h22a == io_addr) begin // @[Ram.scala 19:35]
          mem_554 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h22b == io_addr) begin // @[Ram.scala 19:35]
          mem_555 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h22c == io_addr) begin // @[Ram.scala 19:35]
          mem_556 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h22d == io_addr) begin // @[Ram.scala 19:35]
          mem_557 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h22e == io_addr) begin // @[Ram.scala 19:35]
          mem_558 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h22f == io_addr) begin // @[Ram.scala 19:35]
          mem_559 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h230 == io_addr) begin // @[Ram.scala 19:35]
          mem_560 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h231 == io_addr) begin // @[Ram.scala 19:35]
          mem_561 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h232 == io_addr) begin // @[Ram.scala 19:35]
          mem_562 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h233 == io_addr) begin // @[Ram.scala 19:35]
          mem_563 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h234 == io_addr) begin // @[Ram.scala 19:35]
          mem_564 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h235 == io_addr) begin // @[Ram.scala 19:35]
          mem_565 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h236 == io_addr) begin // @[Ram.scala 19:35]
          mem_566 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h237 == io_addr) begin // @[Ram.scala 19:35]
          mem_567 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h238 == io_addr) begin // @[Ram.scala 19:35]
          mem_568 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h239 == io_addr) begin // @[Ram.scala 19:35]
          mem_569 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h23a == io_addr) begin // @[Ram.scala 19:35]
          mem_570 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h23b == io_addr) begin // @[Ram.scala 19:35]
          mem_571 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h23c == io_addr) begin // @[Ram.scala 19:35]
          mem_572 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h23d == io_addr) begin // @[Ram.scala 19:35]
          mem_573 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h23e == io_addr) begin // @[Ram.scala 19:35]
          mem_574 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h23f == io_addr) begin // @[Ram.scala 19:35]
          mem_575 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h240 == io_addr) begin // @[Ram.scala 19:35]
          mem_576 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h241 == io_addr) begin // @[Ram.scala 19:35]
          mem_577 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h242 == io_addr) begin // @[Ram.scala 19:35]
          mem_578 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h243 == io_addr) begin // @[Ram.scala 19:35]
          mem_579 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h244 == io_addr) begin // @[Ram.scala 19:35]
          mem_580 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h245 == io_addr) begin // @[Ram.scala 19:35]
          mem_581 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h246 == io_addr) begin // @[Ram.scala 19:35]
          mem_582 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h247 == io_addr) begin // @[Ram.scala 19:35]
          mem_583 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h248 == io_addr) begin // @[Ram.scala 19:35]
          mem_584 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h249 == io_addr) begin // @[Ram.scala 19:35]
          mem_585 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h24a == io_addr) begin // @[Ram.scala 19:35]
          mem_586 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h24b == io_addr) begin // @[Ram.scala 19:35]
          mem_587 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h24c == io_addr) begin // @[Ram.scala 19:35]
          mem_588 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h24d == io_addr) begin // @[Ram.scala 19:35]
          mem_589 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h24e == io_addr) begin // @[Ram.scala 19:35]
          mem_590 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h24f == io_addr) begin // @[Ram.scala 19:35]
          mem_591 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h250 == io_addr) begin // @[Ram.scala 19:35]
          mem_592 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h251 == io_addr) begin // @[Ram.scala 19:35]
          mem_593 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h252 == io_addr) begin // @[Ram.scala 19:35]
          mem_594 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h253 == io_addr) begin // @[Ram.scala 19:35]
          mem_595 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h254 == io_addr) begin // @[Ram.scala 19:35]
          mem_596 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h255 == io_addr) begin // @[Ram.scala 19:35]
          mem_597 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h256 == io_addr) begin // @[Ram.scala 19:35]
          mem_598 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h257 == io_addr) begin // @[Ram.scala 19:35]
          mem_599 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h258 == io_addr) begin // @[Ram.scala 19:35]
          mem_600 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h259 == io_addr) begin // @[Ram.scala 19:35]
          mem_601 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h25a == io_addr) begin // @[Ram.scala 19:35]
          mem_602 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h25b == io_addr) begin // @[Ram.scala 19:35]
          mem_603 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h25c == io_addr) begin // @[Ram.scala 19:35]
          mem_604 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h25d == io_addr) begin // @[Ram.scala 19:35]
          mem_605 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h25e == io_addr) begin // @[Ram.scala 19:35]
          mem_606 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h25f == io_addr) begin // @[Ram.scala 19:35]
          mem_607 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h260 == io_addr) begin // @[Ram.scala 19:35]
          mem_608 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h261 == io_addr) begin // @[Ram.scala 19:35]
          mem_609 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h262 == io_addr) begin // @[Ram.scala 19:35]
          mem_610 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h263 == io_addr) begin // @[Ram.scala 19:35]
          mem_611 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h264 == io_addr) begin // @[Ram.scala 19:35]
          mem_612 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h265 == io_addr) begin // @[Ram.scala 19:35]
          mem_613 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h266 == io_addr) begin // @[Ram.scala 19:35]
          mem_614 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h267 == io_addr) begin // @[Ram.scala 19:35]
          mem_615 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h268 == io_addr) begin // @[Ram.scala 19:35]
          mem_616 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h269 == io_addr) begin // @[Ram.scala 19:35]
          mem_617 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h26a == io_addr) begin // @[Ram.scala 19:35]
          mem_618 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h26b == io_addr) begin // @[Ram.scala 19:35]
          mem_619 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h26c == io_addr) begin // @[Ram.scala 19:35]
          mem_620 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h26d == io_addr) begin // @[Ram.scala 19:35]
          mem_621 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h26e == io_addr) begin // @[Ram.scala 19:35]
          mem_622 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h26f == io_addr) begin // @[Ram.scala 19:35]
          mem_623 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h270 == io_addr) begin // @[Ram.scala 19:35]
          mem_624 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h271 == io_addr) begin // @[Ram.scala 19:35]
          mem_625 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h272 == io_addr) begin // @[Ram.scala 19:35]
          mem_626 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h273 == io_addr) begin // @[Ram.scala 19:35]
          mem_627 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h274 == io_addr) begin // @[Ram.scala 19:35]
          mem_628 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h275 == io_addr) begin // @[Ram.scala 19:35]
          mem_629 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h276 == io_addr) begin // @[Ram.scala 19:35]
          mem_630 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h277 == io_addr) begin // @[Ram.scala 19:35]
          mem_631 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h278 == io_addr) begin // @[Ram.scala 19:35]
          mem_632 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h279 == io_addr) begin // @[Ram.scala 19:35]
          mem_633 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h27a == io_addr) begin // @[Ram.scala 19:35]
          mem_634 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h27b == io_addr) begin // @[Ram.scala 19:35]
          mem_635 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h27c == io_addr) begin // @[Ram.scala 19:35]
          mem_636 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h27d == io_addr) begin // @[Ram.scala 19:35]
          mem_637 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h27e == io_addr) begin // @[Ram.scala 19:35]
          mem_638 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h27f == io_addr) begin // @[Ram.scala 19:35]
          mem_639 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h280 == io_addr) begin // @[Ram.scala 19:35]
          mem_640 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h281 == io_addr) begin // @[Ram.scala 19:35]
          mem_641 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h282 == io_addr) begin // @[Ram.scala 19:35]
          mem_642 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h283 == io_addr) begin // @[Ram.scala 19:35]
          mem_643 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h284 == io_addr) begin // @[Ram.scala 19:35]
          mem_644 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h285 == io_addr) begin // @[Ram.scala 19:35]
          mem_645 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h286 == io_addr) begin // @[Ram.scala 19:35]
          mem_646 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h287 == io_addr) begin // @[Ram.scala 19:35]
          mem_647 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h288 == io_addr) begin // @[Ram.scala 19:35]
          mem_648 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h289 == io_addr) begin // @[Ram.scala 19:35]
          mem_649 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h28a == io_addr) begin // @[Ram.scala 19:35]
          mem_650 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h28b == io_addr) begin // @[Ram.scala 19:35]
          mem_651 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h28c == io_addr) begin // @[Ram.scala 19:35]
          mem_652 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h28d == io_addr) begin // @[Ram.scala 19:35]
          mem_653 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h28e == io_addr) begin // @[Ram.scala 19:35]
          mem_654 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h28f == io_addr) begin // @[Ram.scala 19:35]
          mem_655 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h290 == io_addr) begin // @[Ram.scala 19:35]
          mem_656 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h291 == io_addr) begin // @[Ram.scala 19:35]
          mem_657 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h292 == io_addr) begin // @[Ram.scala 19:35]
          mem_658 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h293 == io_addr) begin // @[Ram.scala 19:35]
          mem_659 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h294 == io_addr) begin // @[Ram.scala 19:35]
          mem_660 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h295 == io_addr) begin // @[Ram.scala 19:35]
          mem_661 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h296 == io_addr) begin // @[Ram.scala 19:35]
          mem_662 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h297 == io_addr) begin // @[Ram.scala 19:35]
          mem_663 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h298 == io_addr) begin // @[Ram.scala 19:35]
          mem_664 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h299 == io_addr) begin // @[Ram.scala 19:35]
          mem_665 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h29a == io_addr) begin // @[Ram.scala 19:35]
          mem_666 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h29b == io_addr) begin // @[Ram.scala 19:35]
          mem_667 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h29c == io_addr) begin // @[Ram.scala 19:35]
          mem_668 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h29d == io_addr) begin // @[Ram.scala 19:35]
          mem_669 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h29e == io_addr) begin // @[Ram.scala 19:35]
          mem_670 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h29f == io_addr) begin // @[Ram.scala 19:35]
          mem_671 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2a0 == io_addr) begin // @[Ram.scala 19:35]
          mem_672 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2a1 == io_addr) begin // @[Ram.scala 19:35]
          mem_673 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2a2 == io_addr) begin // @[Ram.scala 19:35]
          mem_674 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2a3 == io_addr) begin // @[Ram.scala 19:35]
          mem_675 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2a4 == io_addr) begin // @[Ram.scala 19:35]
          mem_676 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2a5 == io_addr) begin // @[Ram.scala 19:35]
          mem_677 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2a6 == io_addr) begin // @[Ram.scala 19:35]
          mem_678 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2a7 == io_addr) begin // @[Ram.scala 19:35]
          mem_679 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2a8 == io_addr) begin // @[Ram.scala 19:35]
          mem_680 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2a9 == io_addr) begin // @[Ram.scala 19:35]
          mem_681 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2aa == io_addr) begin // @[Ram.scala 19:35]
          mem_682 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ab == io_addr) begin // @[Ram.scala 19:35]
          mem_683 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ac == io_addr) begin // @[Ram.scala 19:35]
          mem_684 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ad == io_addr) begin // @[Ram.scala 19:35]
          mem_685 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ae == io_addr) begin // @[Ram.scala 19:35]
          mem_686 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2af == io_addr) begin // @[Ram.scala 19:35]
          mem_687 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2b0 == io_addr) begin // @[Ram.scala 19:35]
          mem_688 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2b1 == io_addr) begin // @[Ram.scala 19:35]
          mem_689 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2b2 == io_addr) begin // @[Ram.scala 19:35]
          mem_690 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2b3 == io_addr) begin // @[Ram.scala 19:35]
          mem_691 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2b4 == io_addr) begin // @[Ram.scala 19:35]
          mem_692 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2b5 == io_addr) begin // @[Ram.scala 19:35]
          mem_693 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2b6 == io_addr) begin // @[Ram.scala 19:35]
          mem_694 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2b7 == io_addr) begin // @[Ram.scala 19:35]
          mem_695 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2b8 == io_addr) begin // @[Ram.scala 19:35]
          mem_696 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2b9 == io_addr) begin // @[Ram.scala 19:35]
          mem_697 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ba == io_addr) begin // @[Ram.scala 19:35]
          mem_698 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2bb == io_addr) begin // @[Ram.scala 19:35]
          mem_699 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2bc == io_addr) begin // @[Ram.scala 19:35]
          mem_700 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2bd == io_addr) begin // @[Ram.scala 19:35]
          mem_701 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2be == io_addr) begin // @[Ram.scala 19:35]
          mem_702 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2bf == io_addr) begin // @[Ram.scala 19:35]
          mem_703 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2c0 == io_addr) begin // @[Ram.scala 19:35]
          mem_704 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2c1 == io_addr) begin // @[Ram.scala 19:35]
          mem_705 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2c2 == io_addr) begin // @[Ram.scala 19:35]
          mem_706 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2c3 == io_addr) begin // @[Ram.scala 19:35]
          mem_707 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2c4 == io_addr) begin // @[Ram.scala 19:35]
          mem_708 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2c5 == io_addr) begin // @[Ram.scala 19:35]
          mem_709 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2c6 == io_addr) begin // @[Ram.scala 19:35]
          mem_710 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2c7 == io_addr) begin // @[Ram.scala 19:35]
          mem_711 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2c8 == io_addr) begin // @[Ram.scala 19:35]
          mem_712 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2c9 == io_addr) begin // @[Ram.scala 19:35]
          mem_713 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ca == io_addr) begin // @[Ram.scala 19:35]
          mem_714 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2cb == io_addr) begin // @[Ram.scala 19:35]
          mem_715 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2cc == io_addr) begin // @[Ram.scala 19:35]
          mem_716 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2cd == io_addr) begin // @[Ram.scala 19:35]
          mem_717 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ce == io_addr) begin // @[Ram.scala 19:35]
          mem_718 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2cf == io_addr) begin // @[Ram.scala 19:35]
          mem_719 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2d0 == io_addr) begin // @[Ram.scala 19:35]
          mem_720 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2d1 == io_addr) begin // @[Ram.scala 19:35]
          mem_721 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2d2 == io_addr) begin // @[Ram.scala 19:35]
          mem_722 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2d3 == io_addr) begin // @[Ram.scala 19:35]
          mem_723 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2d4 == io_addr) begin // @[Ram.scala 19:35]
          mem_724 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2d5 == io_addr) begin // @[Ram.scala 19:35]
          mem_725 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2d6 == io_addr) begin // @[Ram.scala 19:35]
          mem_726 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2d7 == io_addr) begin // @[Ram.scala 19:35]
          mem_727 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2d8 == io_addr) begin // @[Ram.scala 19:35]
          mem_728 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2d9 == io_addr) begin // @[Ram.scala 19:35]
          mem_729 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2da == io_addr) begin // @[Ram.scala 19:35]
          mem_730 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2db == io_addr) begin // @[Ram.scala 19:35]
          mem_731 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2dc == io_addr) begin // @[Ram.scala 19:35]
          mem_732 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2dd == io_addr) begin // @[Ram.scala 19:35]
          mem_733 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2de == io_addr) begin // @[Ram.scala 19:35]
          mem_734 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2df == io_addr) begin // @[Ram.scala 19:35]
          mem_735 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2e0 == io_addr) begin // @[Ram.scala 19:35]
          mem_736 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2e1 == io_addr) begin // @[Ram.scala 19:35]
          mem_737 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2e2 == io_addr) begin // @[Ram.scala 19:35]
          mem_738 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2e3 == io_addr) begin // @[Ram.scala 19:35]
          mem_739 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2e4 == io_addr) begin // @[Ram.scala 19:35]
          mem_740 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2e5 == io_addr) begin // @[Ram.scala 19:35]
          mem_741 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2e6 == io_addr) begin // @[Ram.scala 19:35]
          mem_742 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2e7 == io_addr) begin // @[Ram.scala 19:35]
          mem_743 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2e8 == io_addr) begin // @[Ram.scala 19:35]
          mem_744 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2e9 == io_addr) begin // @[Ram.scala 19:35]
          mem_745 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ea == io_addr) begin // @[Ram.scala 19:35]
          mem_746 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2eb == io_addr) begin // @[Ram.scala 19:35]
          mem_747 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ec == io_addr) begin // @[Ram.scala 19:35]
          mem_748 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ed == io_addr) begin // @[Ram.scala 19:35]
          mem_749 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ee == io_addr) begin // @[Ram.scala 19:35]
          mem_750 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ef == io_addr) begin // @[Ram.scala 19:35]
          mem_751 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2f0 == io_addr) begin // @[Ram.scala 19:35]
          mem_752 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2f1 == io_addr) begin // @[Ram.scala 19:35]
          mem_753 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2f2 == io_addr) begin // @[Ram.scala 19:35]
          mem_754 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2f3 == io_addr) begin // @[Ram.scala 19:35]
          mem_755 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2f4 == io_addr) begin // @[Ram.scala 19:35]
          mem_756 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2f5 == io_addr) begin // @[Ram.scala 19:35]
          mem_757 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2f6 == io_addr) begin // @[Ram.scala 19:35]
          mem_758 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2f7 == io_addr) begin // @[Ram.scala 19:35]
          mem_759 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2f8 == io_addr) begin // @[Ram.scala 19:35]
          mem_760 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2f9 == io_addr) begin // @[Ram.scala 19:35]
          mem_761 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2fa == io_addr) begin // @[Ram.scala 19:35]
          mem_762 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2fb == io_addr) begin // @[Ram.scala 19:35]
          mem_763 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2fc == io_addr) begin // @[Ram.scala 19:35]
          mem_764 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2fd == io_addr) begin // @[Ram.scala 19:35]
          mem_765 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2fe == io_addr) begin // @[Ram.scala 19:35]
          mem_766 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h2ff == io_addr) begin // @[Ram.scala 19:35]
          mem_767 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h300 == io_addr) begin // @[Ram.scala 19:35]
          mem_768 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h301 == io_addr) begin // @[Ram.scala 19:35]
          mem_769 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h302 == io_addr) begin // @[Ram.scala 19:35]
          mem_770 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h303 == io_addr) begin // @[Ram.scala 19:35]
          mem_771 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h304 == io_addr) begin // @[Ram.scala 19:35]
          mem_772 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h305 == io_addr) begin // @[Ram.scala 19:35]
          mem_773 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h306 == io_addr) begin // @[Ram.scala 19:35]
          mem_774 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h307 == io_addr) begin // @[Ram.scala 19:35]
          mem_775 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h308 == io_addr) begin // @[Ram.scala 19:35]
          mem_776 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h309 == io_addr) begin // @[Ram.scala 19:35]
          mem_777 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h30a == io_addr) begin // @[Ram.scala 19:35]
          mem_778 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h30b == io_addr) begin // @[Ram.scala 19:35]
          mem_779 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h30c == io_addr) begin // @[Ram.scala 19:35]
          mem_780 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h30d == io_addr) begin // @[Ram.scala 19:35]
          mem_781 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h30e == io_addr) begin // @[Ram.scala 19:35]
          mem_782 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h30f == io_addr) begin // @[Ram.scala 19:35]
          mem_783 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h310 == io_addr) begin // @[Ram.scala 19:35]
          mem_784 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h311 == io_addr) begin // @[Ram.scala 19:35]
          mem_785 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h312 == io_addr) begin // @[Ram.scala 19:35]
          mem_786 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h313 == io_addr) begin // @[Ram.scala 19:35]
          mem_787 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h314 == io_addr) begin // @[Ram.scala 19:35]
          mem_788 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h315 == io_addr) begin // @[Ram.scala 19:35]
          mem_789 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h316 == io_addr) begin // @[Ram.scala 19:35]
          mem_790 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h317 == io_addr) begin // @[Ram.scala 19:35]
          mem_791 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h318 == io_addr) begin // @[Ram.scala 19:35]
          mem_792 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h319 == io_addr) begin // @[Ram.scala 19:35]
          mem_793 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h31a == io_addr) begin // @[Ram.scala 19:35]
          mem_794 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h31b == io_addr) begin // @[Ram.scala 19:35]
          mem_795 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h31c == io_addr) begin // @[Ram.scala 19:35]
          mem_796 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h31d == io_addr) begin // @[Ram.scala 19:35]
          mem_797 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h31e == io_addr) begin // @[Ram.scala 19:35]
          mem_798 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h31f == io_addr) begin // @[Ram.scala 19:35]
          mem_799 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h320 == io_addr) begin // @[Ram.scala 19:35]
          mem_800 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h321 == io_addr) begin // @[Ram.scala 19:35]
          mem_801 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h322 == io_addr) begin // @[Ram.scala 19:35]
          mem_802 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h323 == io_addr) begin // @[Ram.scala 19:35]
          mem_803 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h324 == io_addr) begin // @[Ram.scala 19:35]
          mem_804 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h325 == io_addr) begin // @[Ram.scala 19:35]
          mem_805 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h326 == io_addr) begin // @[Ram.scala 19:35]
          mem_806 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h327 == io_addr) begin // @[Ram.scala 19:35]
          mem_807 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h328 == io_addr) begin // @[Ram.scala 19:35]
          mem_808 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h329 == io_addr) begin // @[Ram.scala 19:35]
          mem_809 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h32a == io_addr) begin // @[Ram.scala 19:35]
          mem_810 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h32b == io_addr) begin // @[Ram.scala 19:35]
          mem_811 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h32c == io_addr) begin // @[Ram.scala 19:35]
          mem_812 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h32d == io_addr) begin // @[Ram.scala 19:35]
          mem_813 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h32e == io_addr) begin // @[Ram.scala 19:35]
          mem_814 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h32f == io_addr) begin // @[Ram.scala 19:35]
          mem_815 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h330 == io_addr) begin // @[Ram.scala 19:35]
          mem_816 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h331 == io_addr) begin // @[Ram.scala 19:35]
          mem_817 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h332 == io_addr) begin // @[Ram.scala 19:35]
          mem_818 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h333 == io_addr) begin // @[Ram.scala 19:35]
          mem_819 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h334 == io_addr) begin // @[Ram.scala 19:35]
          mem_820 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h335 == io_addr) begin // @[Ram.scala 19:35]
          mem_821 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h336 == io_addr) begin // @[Ram.scala 19:35]
          mem_822 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h337 == io_addr) begin // @[Ram.scala 19:35]
          mem_823 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h338 == io_addr) begin // @[Ram.scala 19:35]
          mem_824 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h339 == io_addr) begin // @[Ram.scala 19:35]
          mem_825 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h33a == io_addr) begin // @[Ram.scala 19:35]
          mem_826 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h33b == io_addr) begin // @[Ram.scala 19:35]
          mem_827 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h33c == io_addr) begin // @[Ram.scala 19:35]
          mem_828 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h33d == io_addr) begin // @[Ram.scala 19:35]
          mem_829 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h33e == io_addr) begin // @[Ram.scala 19:35]
          mem_830 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h33f == io_addr) begin // @[Ram.scala 19:35]
          mem_831 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h340 == io_addr) begin // @[Ram.scala 19:35]
          mem_832 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h341 == io_addr) begin // @[Ram.scala 19:35]
          mem_833 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h342 == io_addr) begin // @[Ram.scala 19:35]
          mem_834 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h343 == io_addr) begin // @[Ram.scala 19:35]
          mem_835 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h344 == io_addr) begin // @[Ram.scala 19:35]
          mem_836 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h345 == io_addr) begin // @[Ram.scala 19:35]
          mem_837 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h346 == io_addr) begin // @[Ram.scala 19:35]
          mem_838 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h347 == io_addr) begin // @[Ram.scala 19:35]
          mem_839 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h348 == io_addr) begin // @[Ram.scala 19:35]
          mem_840 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h349 == io_addr) begin // @[Ram.scala 19:35]
          mem_841 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h34a == io_addr) begin // @[Ram.scala 19:35]
          mem_842 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h34b == io_addr) begin // @[Ram.scala 19:35]
          mem_843 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h34c == io_addr) begin // @[Ram.scala 19:35]
          mem_844 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h34d == io_addr) begin // @[Ram.scala 19:35]
          mem_845 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h34e == io_addr) begin // @[Ram.scala 19:35]
          mem_846 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h34f == io_addr) begin // @[Ram.scala 19:35]
          mem_847 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h350 == io_addr) begin // @[Ram.scala 19:35]
          mem_848 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h351 == io_addr) begin // @[Ram.scala 19:35]
          mem_849 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h352 == io_addr) begin // @[Ram.scala 19:35]
          mem_850 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h353 == io_addr) begin // @[Ram.scala 19:35]
          mem_851 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h354 == io_addr) begin // @[Ram.scala 19:35]
          mem_852 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h355 == io_addr) begin // @[Ram.scala 19:35]
          mem_853 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h356 == io_addr) begin // @[Ram.scala 19:35]
          mem_854 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h357 == io_addr) begin // @[Ram.scala 19:35]
          mem_855 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h358 == io_addr) begin // @[Ram.scala 19:35]
          mem_856 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h359 == io_addr) begin // @[Ram.scala 19:35]
          mem_857 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h35a == io_addr) begin // @[Ram.scala 19:35]
          mem_858 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h35b == io_addr) begin // @[Ram.scala 19:35]
          mem_859 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h35c == io_addr) begin // @[Ram.scala 19:35]
          mem_860 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h35d == io_addr) begin // @[Ram.scala 19:35]
          mem_861 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h35e == io_addr) begin // @[Ram.scala 19:35]
          mem_862 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h35f == io_addr) begin // @[Ram.scala 19:35]
          mem_863 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h360 == io_addr) begin // @[Ram.scala 19:35]
          mem_864 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h361 == io_addr) begin // @[Ram.scala 19:35]
          mem_865 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h362 == io_addr) begin // @[Ram.scala 19:35]
          mem_866 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h363 == io_addr) begin // @[Ram.scala 19:35]
          mem_867 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h364 == io_addr) begin // @[Ram.scala 19:35]
          mem_868 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h365 == io_addr) begin // @[Ram.scala 19:35]
          mem_869 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h366 == io_addr) begin // @[Ram.scala 19:35]
          mem_870 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h367 == io_addr) begin // @[Ram.scala 19:35]
          mem_871 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h368 == io_addr) begin // @[Ram.scala 19:35]
          mem_872 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h369 == io_addr) begin // @[Ram.scala 19:35]
          mem_873 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h36a == io_addr) begin // @[Ram.scala 19:35]
          mem_874 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h36b == io_addr) begin // @[Ram.scala 19:35]
          mem_875 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h36c == io_addr) begin // @[Ram.scala 19:35]
          mem_876 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h36d == io_addr) begin // @[Ram.scala 19:35]
          mem_877 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h36e == io_addr) begin // @[Ram.scala 19:35]
          mem_878 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h36f == io_addr) begin // @[Ram.scala 19:35]
          mem_879 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h370 == io_addr) begin // @[Ram.scala 19:35]
          mem_880 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h371 == io_addr) begin // @[Ram.scala 19:35]
          mem_881 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h372 == io_addr) begin // @[Ram.scala 19:35]
          mem_882 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h373 == io_addr) begin // @[Ram.scala 19:35]
          mem_883 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h374 == io_addr) begin // @[Ram.scala 19:35]
          mem_884 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h375 == io_addr) begin // @[Ram.scala 19:35]
          mem_885 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h376 == io_addr) begin // @[Ram.scala 19:35]
          mem_886 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h377 == io_addr) begin // @[Ram.scala 19:35]
          mem_887 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h378 == io_addr) begin // @[Ram.scala 19:35]
          mem_888 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h379 == io_addr) begin // @[Ram.scala 19:35]
          mem_889 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h37a == io_addr) begin // @[Ram.scala 19:35]
          mem_890 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h37b == io_addr) begin // @[Ram.scala 19:35]
          mem_891 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h37c == io_addr) begin // @[Ram.scala 19:35]
          mem_892 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h37d == io_addr) begin // @[Ram.scala 19:35]
          mem_893 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h37e == io_addr) begin // @[Ram.scala 19:35]
          mem_894 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h37f == io_addr) begin // @[Ram.scala 19:35]
          mem_895 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h380 == io_addr) begin // @[Ram.scala 19:35]
          mem_896 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h381 == io_addr) begin // @[Ram.scala 19:35]
          mem_897 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h382 == io_addr) begin // @[Ram.scala 19:35]
          mem_898 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h383 == io_addr) begin // @[Ram.scala 19:35]
          mem_899 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h384 == io_addr) begin // @[Ram.scala 19:35]
          mem_900 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h385 == io_addr) begin // @[Ram.scala 19:35]
          mem_901 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h386 == io_addr) begin // @[Ram.scala 19:35]
          mem_902 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h387 == io_addr) begin // @[Ram.scala 19:35]
          mem_903 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h388 == io_addr) begin // @[Ram.scala 19:35]
          mem_904 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h389 == io_addr) begin // @[Ram.scala 19:35]
          mem_905 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h38a == io_addr) begin // @[Ram.scala 19:35]
          mem_906 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h38b == io_addr) begin // @[Ram.scala 19:35]
          mem_907 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h38c == io_addr) begin // @[Ram.scala 19:35]
          mem_908 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h38d == io_addr) begin // @[Ram.scala 19:35]
          mem_909 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h38e == io_addr) begin // @[Ram.scala 19:35]
          mem_910 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h38f == io_addr) begin // @[Ram.scala 19:35]
          mem_911 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h390 == io_addr) begin // @[Ram.scala 19:35]
          mem_912 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h391 == io_addr) begin // @[Ram.scala 19:35]
          mem_913 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h392 == io_addr) begin // @[Ram.scala 19:35]
          mem_914 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h393 == io_addr) begin // @[Ram.scala 19:35]
          mem_915 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h394 == io_addr) begin // @[Ram.scala 19:35]
          mem_916 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h395 == io_addr) begin // @[Ram.scala 19:35]
          mem_917 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h396 == io_addr) begin // @[Ram.scala 19:35]
          mem_918 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h397 == io_addr) begin // @[Ram.scala 19:35]
          mem_919 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h398 == io_addr) begin // @[Ram.scala 19:35]
          mem_920 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h399 == io_addr) begin // @[Ram.scala 19:35]
          mem_921 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h39a == io_addr) begin // @[Ram.scala 19:35]
          mem_922 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h39b == io_addr) begin // @[Ram.scala 19:35]
          mem_923 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h39c == io_addr) begin // @[Ram.scala 19:35]
          mem_924 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h39d == io_addr) begin // @[Ram.scala 19:35]
          mem_925 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h39e == io_addr) begin // @[Ram.scala 19:35]
          mem_926 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h39f == io_addr) begin // @[Ram.scala 19:35]
          mem_927 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3a0 == io_addr) begin // @[Ram.scala 19:35]
          mem_928 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3a1 == io_addr) begin // @[Ram.scala 19:35]
          mem_929 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3a2 == io_addr) begin // @[Ram.scala 19:35]
          mem_930 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3a3 == io_addr) begin // @[Ram.scala 19:35]
          mem_931 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3a4 == io_addr) begin // @[Ram.scala 19:35]
          mem_932 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3a5 == io_addr) begin // @[Ram.scala 19:35]
          mem_933 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3a6 == io_addr) begin // @[Ram.scala 19:35]
          mem_934 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3a7 == io_addr) begin // @[Ram.scala 19:35]
          mem_935 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3a8 == io_addr) begin // @[Ram.scala 19:35]
          mem_936 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3a9 == io_addr) begin // @[Ram.scala 19:35]
          mem_937 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3aa == io_addr) begin // @[Ram.scala 19:35]
          mem_938 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ab == io_addr) begin // @[Ram.scala 19:35]
          mem_939 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ac == io_addr) begin // @[Ram.scala 19:35]
          mem_940 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ad == io_addr) begin // @[Ram.scala 19:35]
          mem_941 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ae == io_addr) begin // @[Ram.scala 19:35]
          mem_942 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3af == io_addr) begin // @[Ram.scala 19:35]
          mem_943 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3b0 == io_addr) begin // @[Ram.scala 19:35]
          mem_944 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3b1 == io_addr) begin // @[Ram.scala 19:35]
          mem_945 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3b2 == io_addr) begin // @[Ram.scala 19:35]
          mem_946 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3b3 == io_addr) begin // @[Ram.scala 19:35]
          mem_947 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3b4 == io_addr) begin // @[Ram.scala 19:35]
          mem_948 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3b5 == io_addr) begin // @[Ram.scala 19:35]
          mem_949 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3b6 == io_addr) begin // @[Ram.scala 19:35]
          mem_950 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3b7 == io_addr) begin // @[Ram.scala 19:35]
          mem_951 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3b8 == io_addr) begin // @[Ram.scala 19:35]
          mem_952 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3b9 == io_addr) begin // @[Ram.scala 19:35]
          mem_953 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ba == io_addr) begin // @[Ram.scala 19:35]
          mem_954 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3bb == io_addr) begin // @[Ram.scala 19:35]
          mem_955 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3bc == io_addr) begin // @[Ram.scala 19:35]
          mem_956 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3bd == io_addr) begin // @[Ram.scala 19:35]
          mem_957 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3be == io_addr) begin // @[Ram.scala 19:35]
          mem_958 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3bf == io_addr) begin // @[Ram.scala 19:35]
          mem_959 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3c0 == io_addr) begin // @[Ram.scala 19:35]
          mem_960 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3c1 == io_addr) begin // @[Ram.scala 19:35]
          mem_961 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3c2 == io_addr) begin // @[Ram.scala 19:35]
          mem_962 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3c3 == io_addr) begin // @[Ram.scala 19:35]
          mem_963 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3c4 == io_addr) begin // @[Ram.scala 19:35]
          mem_964 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3c5 == io_addr) begin // @[Ram.scala 19:35]
          mem_965 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3c6 == io_addr) begin // @[Ram.scala 19:35]
          mem_966 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3c7 == io_addr) begin // @[Ram.scala 19:35]
          mem_967 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3c8 == io_addr) begin // @[Ram.scala 19:35]
          mem_968 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3c9 == io_addr) begin // @[Ram.scala 19:35]
          mem_969 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ca == io_addr) begin // @[Ram.scala 19:35]
          mem_970 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3cb == io_addr) begin // @[Ram.scala 19:35]
          mem_971 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3cc == io_addr) begin // @[Ram.scala 19:35]
          mem_972 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3cd == io_addr) begin // @[Ram.scala 19:35]
          mem_973 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ce == io_addr) begin // @[Ram.scala 19:35]
          mem_974 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3cf == io_addr) begin // @[Ram.scala 19:35]
          mem_975 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3d0 == io_addr) begin // @[Ram.scala 19:35]
          mem_976 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3d1 == io_addr) begin // @[Ram.scala 19:35]
          mem_977 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3d2 == io_addr) begin // @[Ram.scala 19:35]
          mem_978 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3d3 == io_addr) begin // @[Ram.scala 19:35]
          mem_979 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3d4 == io_addr) begin // @[Ram.scala 19:35]
          mem_980 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3d5 == io_addr) begin // @[Ram.scala 19:35]
          mem_981 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3d6 == io_addr) begin // @[Ram.scala 19:35]
          mem_982 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3d7 == io_addr) begin // @[Ram.scala 19:35]
          mem_983 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3d8 == io_addr) begin // @[Ram.scala 19:35]
          mem_984 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3d9 == io_addr) begin // @[Ram.scala 19:35]
          mem_985 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3da == io_addr) begin // @[Ram.scala 19:35]
          mem_986 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3db == io_addr) begin // @[Ram.scala 19:35]
          mem_987 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3dc == io_addr) begin // @[Ram.scala 19:35]
          mem_988 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3dd == io_addr) begin // @[Ram.scala 19:35]
          mem_989 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3de == io_addr) begin // @[Ram.scala 19:35]
          mem_990 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3df == io_addr) begin // @[Ram.scala 19:35]
          mem_991 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3e0 == io_addr) begin // @[Ram.scala 19:35]
          mem_992 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3e1 == io_addr) begin // @[Ram.scala 19:35]
          mem_993 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3e2 == io_addr) begin // @[Ram.scala 19:35]
          mem_994 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3e3 == io_addr) begin // @[Ram.scala 19:35]
          mem_995 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3e4 == io_addr) begin // @[Ram.scala 19:35]
          mem_996 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3e5 == io_addr) begin // @[Ram.scala 19:35]
          mem_997 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3e6 == io_addr) begin // @[Ram.scala 19:35]
          mem_998 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3e7 == io_addr) begin // @[Ram.scala 19:35]
          mem_999 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3e8 == io_addr) begin // @[Ram.scala 19:35]
          mem_1000 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3e9 == io_addr) begin // @[Ram.scala 19:35]
          mem_1001 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ea == io_addr) begin // @[Ram.scala 19:35]
          mem_1002 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3eb == io_addr) begin // @[Ram.scala 19:35]
          mem_1003 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ec == io_addr) begin // @[Ram.scala 19:35]
          mem_1004 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ed == io_addr) begin // @[Ram.scala 19:35]
          mem_1005 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ee == io_addr) begin // @[Ram.scala 19:35]
          mem_1006 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ef == io_addr) begin // @[Ram.scala 19:35]
          mem_1007 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3f0 == io_addr) begin // @[Ram.scala 19:35]
          mem_1008 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3f1 == io_addr) begin // @[Ram.scala 19:35]
          mem_1009 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3f2 == io_addr) begin // @[Ram.scala 19:35]
          mem_1010 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3f3 == io_addr) begin // @[Ram.scala 19:35]
          mem_1011 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3f4 == io_addr) begin // @[Ram.scala 19:35]
          mem_1012 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3f5 == io_addr) begin // @[Ram.scala 19:35]
          mem_1013 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3f6 == io_addr) begin // @[Ram.scala 19:35]
          mem_1014 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3f7 == io_addr) begin // @[Ram.scala 19:35]
          mem_1015 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3f8 == io_addr) begin // @[Ram.scala 19:35]
          mem_1016 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3f9 == io_addr) begin // @[Ram.scala 19:35]
          mem_1017 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3fa == io_addr) begin // @[Ram.scala 19:35]
          mem_1018 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3fb == io_addr) begin // @[Ram.scala 19:35]
          mem_1019 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3fc == io_addr) begin // @[Ram.scala 19:35]
          mem_1020 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3fd == io_addr) begin // @[Ram.scala 19:35]
          mem_1021 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3fe == io_addr) begin // @[Ram.scala 19:35]
          mem_1022 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
    if (io_enable) begin // @[Ram.scala 18:19]
      if (io_write) begin // @[Ram.scala 19:20]
        if (10'h3ff == io_addr) begin // @[Ram.scala 19:35]
          mem_1023 <= io_dataIn; // @[Ram.scala 19:35]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  mem_0 = _RAND_0[255:0];
  _RAND_1 = {8{`RANDOM}};
  mem_1 = _RAND_1[255:0];
  _RAND_2 = {8{`RANDOM}};
  mem_2 = _RAND_2[255:0];
  _RAND_3 = {8{`RANDOM}};
  mem_3 = _RAND_3[255:0];
  _RAND_4 = {8{`RANDOM}};
  mem_4 = _RAND_4[255:0];
  _RAND_5 = {8{`RANDOM}};
  mem_5 = _RAND_5[255:0];
  _RAND_6 = {8{`RANDOM}};
  mem_6 = _RAND_6[255:0];
  _RAND_7 = {8{`RANDOM}};
  mem_7 = _RAND_7[255:0];
  _RAND_8 = {8{`RANDOM}};
  mem_8 = _RAND_8[255:0];
  _RAND_9 = {8{`RANDOM}};
  mem_9 = _RAND_9[255:0];
  _RAND_10 = {8{`RANDOM}};
  mem_10 = _RAND_10[255:0];
  _RAND_11 = {8{`RANDOM}};
  mem_11 = _RAND_11[255:0];
  _RAND_12 = {8{`RANDOM}};
  mem_12 = _RAND_12[255:0];
  _RAND_13 = {8{`RANDOM}};
  mem_13 = _RAND_13[255:0];
  _RAND_14 = {8{`RANDOM}};
  mem_14 = _RAND_14[255:0];
  _RAND_15 = {8{`RANDOM}};
  mem_15 = _RAND_15[255:0];
  _RAND_16 = {8{`RANDOM}};
  mem_16 = _RAND_16[255:0];
  _RAND_17 = {8{`RANDOM}};
  mem_17 = _RAND_17[255:0];
  _RAND_18 = {8{`RANDOM}};
  mem_18 = _RAND_18[255:0];
  _RAND_19 = {8{`RANDOM}};
  mem_19 = _RAND_19[255:0];
  _RAND_20 = {8{`RANDOM}};
  mem_20 = _RAND_20[255:0];
  _RAND_21 = {8{`RANDOM}};
  mem_21 = _RAND_21[255:0];
  _RAND_22 = {8{`RANDOM}};
  mem_22 = _RAND_22[255:0];
  _RAND_23 = {8{`RANDOM}};
  mem_23 = _RAND_23[255:0];
  _RAND_24 = {8{`RANDOM}};
  mem_24 = _RAND_24[255:0];
  _RAND_25 = {8{`RANDOM}};
  mem_25 = _RAND_25[255:0];
  _RAND_26 = {8{`RANDOM}};
  mem_26 = _RAND_26[255:0];
  _RAND_27 = {8{`RANDOM}};
  mem_27 = _RAND_27[255:0];
  _RAND_28 = {8{`RANDOM}};
  mem_28 = _RAND_28[255:0];
  _RAND_29 = {8{`RANDOM}};
  mem_29 = _RAND_29[255:0];
  _RAND_30 = {8{`RANDOM}};
  mem_30 = _RAND_30[255:0];
  _RAND_31 = {8{`RANDOM}};
  mem_31 = _RAND_31[255:0];
  _RAND_32 = {8{`RANDOM}};
  mem_32 = _RAND_32[255:0];
  _RAND_33 = {8{`RANDOM}};
  mem_33 = _RAND_33[255:0];
  _RAND_34 = {8{`RANDOM}};
  mem_34 = _RAND_34[255:0];
  _RAND_35 = {8{`RANDOM}};
  mem_35 = _RAND_35[255:0];
  _RAND_36 = {8{`RANDOM}};
  mem_36 = _RAND_36[255:0];
  _RAND_37 = {8{`RANDOM}};
  mem_37 = _RAND_37[255:0];
  _RAND_38 = {8{`RANDOM}};
  mem_38 = _RAND_38[255:0];
  _RAND_39 = {8{`RANDOM}};
  mem_39 = _RAND_39[255:0];
  _RAND_40 = {8{`RANDOM}};
  mem_40 = _RAND_40[255:0];
  _RAND_41 = {8{`RANDOM}};
  mem_41 = _RAND_41[255:0];
  _RAND_42 = {8{`RANDOM}};
  mem_42 = _RAND_42[255:0];
  _RAND_43 = {8{`RANDOM}};
  mem_43 = _RAND_43[255:0];
  _RAND_44 = {8{`RANDOM}};
  mem_44 = _RAND_44[255:0];
  _RAND_45 = {8{`RANDOM}};
  mem_45 = _RAND_45[255:0];
  _RAND_46 = {8{`RANDOM}};
  mem_46 = _RAND_46[255:0];
  _RAND_47 = {8{`RANDOM}};
  mem_47 = _RAND_47[255:0];
  _RAND_48 = {8{`RANDOM}};
  mem_48 = _RAND_48[255:0];
  _RAND_49 = {8{`RANDOM}};
  mem_49 = _RAND_49[255:0];
  _RAND_50 = {8{`RANDOM}};
  mem_50 = _RAND_50[255:0];
  _RAND_51 = {8{`RANDOM}};
  mem_51 = _RAND_51[255:0];
  _RAND_52 = {8{`RANDOM}};
  mem_52 = _RAND_52[255:0];
  _RAND_53 = {8{`RANDOM}};
  mem_53 = _RAND_53[255:0];
  _RAND_54 = {8{`RANDOM}};
  mem_54 = _RAND_54[255:0];
  _RAND_55 = {8{`RANDOM}};
  mem_55 = _RAND_55[255:0];
  _RAND_56 = {8{`RANDOM}};
  mem_56 = _RAND_56[255:0];
  _RAND_57 = {8{`RANDOM}};
  mem_57 = _RAND_57[255:0];
  _RAND_58 = {8{`RANDOM}};
  mem_58 = _RAND_58[255:0];
  _RAND_59 = {8{`RANDOM}};
  mem_59 = _RAND_59[255:0];
  _RAND_60 = {8{`RANDOM}};
  mem_60 = _RAND_60[255:0];
  _RAND_61 = {8{`RANDOM}};
  mem_61 = _RAND_61[255:0];
  _RAND_62 = {8{`RANDOM}};
  mem_62 = _RAND_62[255:0];
  _RAND_63 = {8{`RANDOM}};
  mem_63 = _RAND_63[255:0];
  _RAND_64 = {8{`RANDOM}};
  mem_64 = _RAND_64[255:0];
  _RAND_65 = {8{`RANDOM}};
  mem_65 = _RAND_65[255:0];
  _RAND_66 = {8{`RANDOM}};
  mem_66 = _RAND_66[255:0];
  _RAND_67 = {8{`RANDOM}};
  mem_67 = _RAND_67[255:0];
  _RAND_68 = {8{`RANDOM}};
  mem_68 = _RAND_68[255:0];
  _RAND_69 = {8{`RANDOM}};
  mem_69 = _RAND_69[255:0];
  _RAND_70 = {8{`RANDOM}};
  mem_70 = _RAND_70[255:0];
  _RAND_71 = {8{`RANDOM}};
  mem_71 = _RAND_71[255:0];
  _RAND_72 = {8{`RANDOM}};
  mem_72 = _RAND_72[255:0];
  _RAND_73 = {8{`RANDOM}};
  mem_73 = _RAND_73[255:0];
  _RAND_74 = {8{`RANDOM}};
  mem_74 = _RAND_74[255:0];
  _RAND_75 = {8{`RANDOM}};
  mem_75 = _RAND_75[255:0];
  _RAND_76 = {8{`RANDOM}};
  mem_76 = _RAND_76[255:0];
  _RAND_77 = {8{`RANDOM}};
  mem_77 = _RAND_77[255:0];
  _RAND_78 = {8{`RANDOM}};
  mem_78 = _RAND_78[255:0];
  _RAND_79 = {8{`RANDOM}};
  mem_79 = _RAND_79[255:0];
  _RAND_80 = {8{`RANDOM}};
  mem_80 = _RAND_80[255:0];
  _RAND_81 = {8{`RANDOM}};
  mem_81 = _RAND_81[255:0];
  _RAND_82 = {8{`RANDOM}};
  mem_82 = _RAND_82[255:0];
  _RAND_83 = {8{`RANDOM}};
  mem_83 = _RAND_83[255:0];
  _RAND_84 = {8{`RANDOM}};
  mem_84 = _RAND_84[255:0];
  _RAND_85 = {8{`RANDOM}};
  mem_85 = _RAND_85[255:0];
  _RAND_86 = {8{`RANDOM}};
  mem_86 = _RAND_86[255:0];
  _RAND_87 = {8{`RANDOM}};
  mem_87 = _RAND_87[255:0];
  _RAND_88 = {8{`RANDOM}};
  mem_88 = _RAND_88[255:0];
  _RAND_89 = {8{`RANDOM}};
  mem_89 = _RAND_89[255:0];
  _RAND_90 = {8{`RANDOM}};
  mem_90 = _RAND_90[255:0];
  _RAND_91 = {8{`RANDOM}};
  mem_91 = _RAND_91[255:0];
  _RAND_92 = {8{`RANDOM}};
  mem_92 = _RAND_92[255:0];
  _RAND_93 = {8{`RANDOM}};
  mem_93 = _RAND_93[255:0];
  _RAND_94 = {8{`RANDOM}};
  mem_94 = _RAND_94[255:0];
  _RAND_95 = {8{`RANDOM}};
  mem_95 = _RAND_95[255:0];
  _RAND_96 = {8{`RANDOM}};
  mem_96 = _RAND_96[255:0];
  _RAND_97 = {8{`RANDOM}};
  mem_97 = _RAND_97[255:0];
  _RAND_98 = {8{`RANDOM}};
  mem_98 = _RAND_98[255:0];
  _RAND_99 = {8{`RANDOM}};
  mem_99 = _RAND_99[255:0];
  _RAND_100 = {8{`RANDOM}};
  mem_100 = _RAND_100[255:0];
  _RAND_101 = {8{`RANDOM}};
  mem_101 = _RAND_101[255:0];
  _RAND_102 = {8{`RANDOM}};
  mem_102 = _RAND_102[255:0];
  _RAND_103 = {8{`RANDOM}};
  mem_103 = _RAND_103[255:0];
  _RAND_104 = {8{`RANDOM}};
  mem_104 = _RAND_104[255:0];
  _RAND_105 = {8{`RANDOM}};
  mem_105 = _RAND_105[255:0];
  _RAND_106 = {8{`RANDOM}};
  mem_106 = _RAND_106[255:0];
  _RAND_107 = {8{`RANDOM}};
  mem_107 = _RAND_107[255:0];
  _RAND_108 = {8{`RANDOM}};
  mem_108 = _RAND_108[255:0];
  _RAND_109 = {8{`RANDOM}};
  mem_109 = _RAND_109[255:0];
  _RAND_110 = {8{`RANDOM}};
  mem_110 = _RAND_110[255:0];
  _RAND_111 = {8{`RANDOM}};
  mem_111 = _RAND_111[255:0];
  _RAND_112 = {8{`RANDOM}};
  mem_112 = _RAND_112[255:0];
  _RAND_113 = {8{`RANDOM}};
  mem_113 = _RAND_113[255:0];
  _RAND_114 = {8{`RANDOM}};
  mem_114 = _RAND_114[255:0];
  _RAND_115 = {8{`RANDOM}};
  mem_115 = _RAND_115[255:0];
  _RAND_116 = {8{`RANDOM}};
  mem_116 = _RAND_116[255:0];
  _RAND_117 = {8{`RANDOM}};
  mem_117 = _RAND_117[255:0];
  _RAND_118 = {8{`RANDOM}};
  mem_118 = _RAND_118[255:0];
  _RAND_119 = {8{`RANDOM}};
  mem_119 = _RAND_119[255:0];
  _RAND_120 = {8{`RANDOM}};
  mem_120 = _RAND_120[255:0];
  _RAND_121 = {8{`RANDOM}};
  mem_121 = _RAND_121[255:0];
  _RAND_122 = {8{`RANDOM}};
  mem_122 = _RAND_122[255:0];
  _RAND_123 = {8{`RANDOM}};
  mem_123 = _RAND_123[255:0];
  _RAND_124 = {8{`RANDOM}};
  mem_124 = _RAND_124[255:0];
  _RAND_125 = {8{`RANDOM}};
  mem_125 = _RAND_125[255:0];
  _RAND_126 = {8{`RANDOM}};
  mem_126 = _RAND_126[255:0];
  _RAND_127 = {8{`RANDOM}};
  mem_127 = _RAND_127[255:0];
  _RAND_128 = {8{`RANDOM}};
  mem_128 = _RAND_128[255:0];
  _RAND_129 = {8{`RANDOM}};
  mem_129 = _RAND_129[255:0];
  _RAND_130 = {8{`RANDOM}};
  mem_130 = _RAND_130[255:0];
  _RAND_131 = {8{`RANDOM}};
  mem_131 = _RAND_131[255:0];
  _RAND_132 = {8{`RANDOM}};
  mem_132 = _RAND_132[255:0];
  _RAND_133 = {8{`RANDOM}};
  mem_133 = _RAND_133[255:0];
  _RAND_134 = {8{`RANDOM}};
  mem_134 = _RAND_134[255:0];
  _RAND_135 = {8{`RANDOM}};
  mem_135 = _RAND_135[255:0];
  _RAND_136 = {8{`RANDOM}};
  mem_136 = _RAND_136[255:0];
  _RAND_137 = {8{`RANDOM}};
  mem_137 = _RAND_137[255:0];
  _RAND_138 = {8{`RANDOM}};
  mem_138 = _RAND_138[255:0];
  _RAND_139 = {8{`RANDOM}};
  mem_139 = _RAND_139[255:0];
  _RAND_140 = {8{`RANDOM}};
  mem_140 = _RAND_140[255:0];
  _RAND_141 = {8{`RANDOM}};
  mem_141 = _RAND_141[255:0];
  _RAND_142 = {8{`RANDOM}};
  mem_142 = _RAND_142[255:0];
  _RAND_143 = {8{`RANDOM}};
  mem_143 = _RAND_143[255:0];
  _RAND_144 = {8{`RANDOM}};
  mem_144 = _RAND_144[255:0];
  _RAND_145 = {8{`RANDOM}};
  mem_145 = _RAND_145[255:0];
  _RAND_146 = {8{`RANDOM}};
  mem_146 = _RAND_146[255:0];
  _RAND_147 = {8{`RANDOM}};
  mem_147 = _RAND_147[255:0];
  _RAND_148 = {8{`RANDOM}};
  mem_148 = _RAND_148[255:0];
  _RAND_149 = {8{`RANDOM}};
  mem_149 = _RAND_149[255:0];
  _RAND_150 = {8{`RANDOM}};
  mem_150 = _RAND_150[255:0];
  _RAND_151 = {8{`RANDOM}};
  mem_151 = _RAND_151[255:0];
  _RAND_152 = {8{`RANDOM}};
  mem_152 = _RAND_152[255:0];
  _RAND_153 = {8{`RANDOM}};
  mem_153 = _RAND_153[255:0];
  _RAND_154 = {8{`RANDOM}};
  mem_154 = _RAND_154[255:0];
  _RAND_155 = {8{`RANDOM}};
  mem_155 = _RAND_155[255:0];
  _RAND_156 = {8{`RANDOM}};
  mem_156 = _RAND_156[255:0];
  _RAND_157 = {8{`RANDOM}};
  mem_157 = _RAND_157[255:0];
  _RAND_158 = {8{`RANDOM}};
  mem_158 = _RAND_158[255:0];
  _RAND_159 = {8{`RANDOM}};
  mem_159 = _RAND_159[255:0];
  _RAND_160 = {8{`RANDOM}};
  mem_160 = _RAND_160[255:0];
  _RAND_161 = {8{`RANDOM}};
  mem_161 = _RAND_161[255:0];
  _RAND_162 = {8{`RANDOM}};
  mem_162 = _RAND_162[255:0];
  _RAND_163 = {8{`RANDOM}};
  mem_163 = _RAND_163[255:0];
  _RAND_164 = {8{`RANDOM}};
  mem_164 = _RAND_164[255:0];
  _RAND_165 = {8{`RANDOM}};
  mem_165 = _RAND_165[255:0];
  _RAND_166 = {8{`RANDOM}};
  mem_166 = _RAND_166[255:0];
  _RAND_167 = {8{`RANDOM}};
  mem_167 = _RAND_167[255:0];
  _RAND_168 = {8{`RANDOM}};
  mem_168 = _RAND_168[255:0];
  _RAND_169 = {8{`RANDOM}};
  mem_169 = _RAND_169[255:0];
  _RAND_170 = {8{`RANDOM}};
  mem_170 = _RAND_170[255:0];
  _RAND_171 = {8{`RANDOM}};
  mem_171 = _RAND_171[255:0];
  _RAND_172 = {8{`RANDOM}};
  mem_172 = _RAND_172[255:0];
  _RAND_173 = {8{`RANDOM}};
  mem_173 = _RAND_173[255:0];
  _RAND_174 = {8{`RANDOM}};
  mem_174 = _RAND_174[255:0];
  _RAND_175 = {8{`RANDOM}};
  mem_175 = _RAND_175[255:0];
  _RAND_176 = {8{`RANDOM}};
  mem_176 = _RAND_176[255:0];
  _RAND_177 = {8{`RANDOM}};
  mem_177 = _RAND_177[255:0];
  _RAND_178 = {8{`RANDOM}};
  mem_178 = _RAND_178[255:0];
  _RAND_179 = {8{`RANDOM}};
  mem_179 = _RAND_179[255:0];
  _RAND_180 = {8{`RANDOM}};
  mem_180 = _RAND_180[255:0];
  _RAND_181 = {8{`RANDOM}};
  mem_181 = _RAND_181[255:0];
  _RAND_182 = {8{`RANDOM}};
  mem_182 = _RAND_182[255:0];
  _RAND_183 = {8{`RANDOM}};
  mem_183 = _RAND_183[255:0];
  _RAND_184 = {8{`RANDOM}};
  mem_184 = _RAND_184[255:0];
  _RAND_185 = {8{`RANDOM}};
  mem_185 = _RAND_185[255:0];
  _RAND_186 = {8{`RANDOM}};
  mem_186 = _RAND_186[255:0];
  _RAND_187 = {8{`RANDOM}};
  mem_187 = _RAND_187[255:0];
  _RAND_188 = {8{`RANDOM}};
  mem_188 = _RAND_188[255:0];
  _RAND_189 = {8{`RANDOM}};
  mem_189 = _RAND_189[255:0];
  _RAND_190 = {8{`RANDOM}};
  mem_190 = _RAND_190[255:0];
  _RAND_191 = {8{`RANDOM}};
  mem_191 = _RAND_191[255:0];
  _RAND_192 = {8{`RANDOM}};
  mem_192 = _RAND_192[255:0];
  _RAND_193 = {8{`RANDOM}};
  mem_193 = _RAND_193[255:0];
  _RAND_194 = {8{`RANDOM}};
  mem_194 = _RAND_194[255:0];
  _RAND_195 = {8{`RANDOM}};
  mem_195 = _RAND_195[255:0];
  _RAND_196 = {8{`RANDOM}};
  mem_196 = _RAND_196[255:0];
  _RAND_197 = {8{`RANDOM}};
  mem_197 = _RAND_197[255:0];
  _RAND_198 = {8{`RANDOM}};
  mem_198 = _RAND_198[255:0];
  _RAND_199 = {8{`RANDOM}};
  mem_199 = _RAND_199[255:0];
  _RAND_200 = {8{`RANDOM}};
  mem_200 = _RAND_200[255:0];
  _RAND_201 = {8{`RANDOM}};
  mem_201 = _RAND_201[255:0];
  _RAND_202 = {8{`RANDOM}};
  mem_202 = _RAND_202[255:0];
  _RAND_203 = {8{`RANDOM}};
  mem_203 = _RAND_203[255:0];
  _RAND_204 = {8{`RANDOM}};
  mem_204 = _RAND_204[255:0];
  _RAND_205 = {8{`RANDOM}};
  mem_205 = _RAND_205[255:0];
  _RAND_206 = {8{`RANDOM}};
  mem_206 = _RAND_206[255:0];
  _RAND_207 = {8{`RANDOM}};
  mem_207 = _RAND_207[255:0];
  _RAND_208 = {8{`RANDOM}};
  mem_208 = _RAND_208[255:0];
  _RAND_209 = {8{`RANDOM}};
  mem_209 = _RAND_209[255:0];
  _RAND_210 = {8{`RANDOM}};
  mem_210 = _RAND_210[255:0];
  _RAND_211 = {8{`RANDOM}};
  mem_211 = _RAND_211[255:0];
  _RAND_212 = {8{`RANDOM}};
  mem_212 = _RAND_212[255:0];
  _RAND_213 = {8{`RANDOM}};
  mem_213 = _RAND_213[255:0];
  _RAND_214 = {8{`RANDOM}};
  mem_214 = _RAND_214[255:0];
  _RAND_215 = {8{`RANDOM}};
  mem_215 = _RAND_215[255:0];
  _RAND_216 = {8{`RANDOM}};
  mem_216 = _RAND_216[255:0];
  _RAND_217 = {8{`RANDOM}};
  mem_217 = _RAND_217[255:0];
  _RAND_218 = {8{`RANDOM}};
  mem_218 = _RAND_218[255:0];
  _RAND_219 = {8{`RANDOM}};
  mem_219 = _RAND_219[255:0];
  _RAND_220 = {8{`RANDOM}};
  mem_220 = _RAND_220[255:0];
  _RAND_221 = {8{`RANDOM}};
  mem_221 = _RAND_221[255:0];
  _RAND_222 = {8{`RANDOM}};
  mem_222 = _RAND_222[255:0];
  _RAND_223 = {8{`RANDOM}};
  mem_223 = _RAND_223[255:0];
  _RAND_224 = {8{`RANDOM}};
  mem_224 = _RAND_224[255:0];
  _RAND_225 = {8{`RANDOM}};
  mem_225 = _RAND_225[255:0];
  _RAND_226 = {8{`RANDOM}};
  mem_226 = _RAND_226[255:0];
  _RAND_227 = {8{`RANDOM}};
  mem_227 = _RAND_227[255:0];
  _RAND_228 = {8{`RANDOM}};
  mem_228 = _RAND_228[255:0];
  _RAND_229 = {8{`RANDOM}};
  mem_229 = _RAND_229[255:0];
  _RAND_230 = {8{`RANDOM}};
  mem_230 = _RAND_230[255:0];
  _RAND_231 = {8{`RANDOM}};
  mem_231 = _RAND_231[255:0];
  _RAND_232 = {8{`RANDOM}};
  mem_232 = _RAND_232[255:0];
  _RAND_233 = {8{`RANDOM}};
  mem_233 = _RAND_233[255:0];
  _RAND_234 = {8{`RANDOM}};
  mem_234 = _RAND_234[255:0];
  _RAND_235 = {8{`RANDOM}};
  mem_235 = _RAND_235[255:0];
  _RAND_236 = {8{`RANDOM}};
  mem_236 = _RAND_236[255:0];
  _RAND_237 = {8{`RANDOM}};
  mem_237 = _RAND_237[255:0];
  _RAND_238 = {8{`RANDOM}};
  mem_238 = _RAND_238[255:0];
  _RAND_239 = {8{`RANDOM}};
  mem_239 = _RAND_239[255:0];
  _RAND_240 = {8{`RANDOM}};
  mem_240 = _RAND_240[255:0];
  _RAND_241 = {8{`RANDOM}};
  mem_241 = _RAND_241[255:0];
  _RAND_242 = {8{`RANDOM}};
  mem_242 = _RAND_242[255:0];
  _RAND_243 = {8{`RANDOM}};
  mem_243 = _RAND_243[255:0];
  _RAND_244 = {8{`RANDOM}};
  mem_244 = _RAND_244[255:0];
  _RAND_245 = {8{`RANDOM}};
  mem_245 = _RAND_245[255:0];
  _RAND_246 = {8{`RANDOM}};
  mem_246 = _RAND_246[255:0];
  _RAND_247 = {8{`RANDOM}};
  mem_247 = _RAND_247[255:0];
  _RAND_248 = {8{`RANDOM}};
  mem_248 = _RAND_248[255:0];
  _RAND_249 = {8{`RANDOM}};
  mem_249 = _RAND_249[255:0];
  _RAND_250 = {8{`RANDOM}};
  mem_250 = _RAND_250[255:0];
  _RAND_251 = {8{`RANDOM}};
  mem_251 = _RAND_251[255:0];
  _RAND_252 = {8{`RANDOM}};
  mem_252 = _RAND_252[255:0];
  _RAND_253 = {8{`RANDOM}};
  mem_253 = _RAND_253[255:0];
  _RAND_254 = {8{`RANDOM}};
  mem_254 = _RAND_254[255:0];
  _RAND_255 = {8{`RANDOM}};
  mem_255 = _RAND_255[255:0];
  _RAND_256 = {8{`RANDOM}};
  mem_256 = _RAND_256[255:0];
  _RAND_257 = {8{`RANDOM}};
  mem_257 = _RAND_257[255:0];
  _RAND_258 = {8{`RANDOM}};
  mem_258 = _RAND_258[255:0];
  _RAND_259 = {8{`RANDOM}};
  mem_259 = _RAND_259[255:0];
  _RAND_260 = {8{`RANDOM}};
  mem_260 = _RAND_260[255:0];
  _RAND_261 = {8{`RANDOM}};
  mem_261 = _RAND_261[255:0];
  _RAND_262 = {8{`RANDOM}};
  mem_262 = _RAND_262[255:0];
  _RAND_263 = {8{`RANDOM}};
  mem_263 = _RAND_263[255:0];
  _RAND_264 = {8{`RANDOM}};
  mem_264 = _RAND_264[255:0];
  _RAND_265 = {8{`RANDOM}};
  mem_265 = _RAND_265[255:0];
  _RAND_266 = {8{`RANDOM}};
  mem_266 = _RAND_266[255:0];
  _RAND_267 = {8{`RANDOM}};
  mem_267 = _RAND_267[255:0];
  _RAND_268 = {8{`RANDOM}};
  mem_268 = _RAND_268[255:0];
  _RAND_269 = {8{`RANDOM}};
  mem_269 = _RAND_269[255:0];
  _RAND_270 = {8{`RANDOM}};
  mem_270 = _RAND_270[255:0];
  _RAND_271 = {8{`RANDOM}};
  mem_271 = _RAND_271[255:0];
  _RAND_272 = {8{`RANDOM}};
  mem_272 = _RAND_272[255:0];
  _RAND_273 = {8{`RANDOM}};
  mem_273 = _RAND_273[255:0];
  _RAND_274 = {8{`RANDOM}};
  mem_274 = _RAND_274[255:0];
  _RAND_275 = {8{`RANDOM}};
  mem_275 = _RAND_275[255:0];
  _RAND_276 = {8{`RANDOM}};
  mem_276 = _RAND_276[255:0];
  _RAND_277 = {8{`RANDOM}};
  mem_277 = _RAND_277[255:0];
  _RAND_278 = {8{`RANDOM}};
  mem_278 = _RAND_278[255:0];
  _RAND_279 = {8{`RANDOM}};
  mem_279 = _RAND_279[255:0];
  _RAND_280 = {8{`RANDOM}};
  mem_280 = _RAND_280[255:0];
  _RAND_281 = {8{`RANDOM}};
  mem_281 = _RAND_281[255:0];
  _RAND_282 = {8{`RANDOM}};
  mem_282 = _RAND_282[255:0];
  _RAND_283 = {8{`RANDOM}};
  mem_283 = _RAND_283[255:0];
  _RAND_284 = {8{`RANDOM}};
  mem_284 = _RAND_284[255:0];
  _RAND_285 = {8{`RANDOM}};
  mem_285 = _RAND_285[255:0];
  _RAND_286 = {8{`RANDOM}};
  mem_286 = _RAND_286[255:0];
  _RAND_287 = {8{`RANDOM}};
  mem_287 = _RAND_287[255:0];
  _RAND_288 = {8{`RANDOM}};
  mem_288 = _RAND_288[255:0];
  _RAND_289 = {8{`RANDOM}};
  mem_289 = _RAND_289[255:0];
  _RAND_290 = {8{`RANDOM}};
  mem_290 = _RAND_290[255:0];
  _RAND_291 = {8{`RANDOM}};
  mem_291 = _RAND_291[255:0];
  _RAND_292 = {8{`RANDOM}};
  mem_292 = _RAND_292[255:0];
  _RAND_293 = {8{`RANDOM}};
  mem_293 = _RAND_293[255:0];
  _RAND_294 = {8{`RANDOM}};
  mem_294 = _RAND_294[255:0];
  _RAND_295 = {8{`RANDOM}};
  mem_295 = _RAND_295[255:0];
  _RAND_296 = {8{`RANDOM}};
  mem_296 = _RAND_296[255:0];
  _RAND_297 = {8{`RANDOM}};
  mem_297 = _RAND_297[255:0];
  _RAND_298 = {8{`RANDOM}};
  mem_298 = _RAND_298[255:0];
  _RAND_299 = {8{`RANDOM}};
  mem_299 = _RAND_299[255:0];
  _RAND_300 = {8{`RANDOM}};
  mem_300 = _RAND_300[255:0];
  _RAND_301 = {8{`RANDOM}};
  mem_301 = _RAND_301[255:0];
  _RAND_302 = {8{`RANDOM}};
  mem_302 = _RAND_302[255:0];
  _RAND_303 = {8{`RANDOM}};
  mem_303 = _RAND_303[255:0];
  _RAND_304 = {8{`RANDOM}};
  mem_304 = _RAND_304[255:0];
  _RAND_305 = {8{`RANDOM}};
  mem_305 = _RAND_305[255:0];
  _RAND_306 = {8{`RANDOM}};
  mem_306 = _RAND_306[255:0];
  _RAND_307 = {8{`RANDOM}};
  mem_307 = _RAND_307[255:0];
  _RAND_308 = {8{`RANDOM}};
  mem_308 = _RAND_308[255:0];
  _RAND_309 = {8{`RANDOM}};
  mem_309 = _RAND_309[255:0];
  _RAND_310 = {8{`RANDOM}};
  mem_310 = _RAND_310[255:0];
  _RAND_311 = {8{`RANDOM}};
  mem_311 = _RAND_311[255:0];
  _RAND_312 = {8{`RANDOM}};
  mem_312 = _RAND_312[255:0];
  _RAND_313 = {8{`RANDOM}};
  mem_313 = _RAND_313[255:0];
  _RAND_314 = {8{`RANDOM}};
  mem_314 = _RAND_314[255:0];
  _RAND_315 = {8{`RANDOM}};
  mem_315 = _RAND_315[255:0];
  _RAND_316 = {8{`RANDOM}};
  mem_316 = _RAND_316[255:0];
  _RAND_317 = {8{`RANDOM}};
  mem_317 = _RAND_317[255:0];
  _RAND_318 = {8{`RANDOM}};
  mem_318 = _RAND_318[255:0];
  _RAND_319 = {8{`RANDOM}};
  mem_319 = _RAND_319[255:0];
  _RAND_320 = {8{`RANDOM}};
  mem_320 = _RAND_320[255:0];
  _RAND_321 = {8{`RANDOM}};
  mem_321 = _RAND_321[255:0];
  _RAND_322 = {8{`RANDOM}};
  mem_322 = _RAND_322[255:0];
  _RAND_323 = {8{`RANDOM}};
  mem_323 = _RAND_323[255:0];
  _RAND_324 = {8{`RANDOM}};
  mem_324 = _RAND_324[255:0];
  _RAND_325 = {8{`RANDOM}};
  mem_325 = _RAND_325[255:0];
  _RAND_326 = {8{`RANDOM}};
  mem_326 = _RAND_326[255:0];
  _RAND_327 = {8{`RANDOM}};
  mem_327 = _RAND_327[255:0];
  _RAND_328 = {8{`RANDOM}};
  mem_328 = _RAND_328[255:0];
  _RAND_329 = {8{`RANDOM}};
  mem_329 = _RAND_329[255:0];
  _RAND_330 = {8{`RANDOM}};
  mem_330 = _RAND_330[255:0];
  _RAND_331 = {8{`RANDOM}};
  mem_331 = _RAND_331[255:0];
  _RAND_332 = {8{`RANDOM}};
  mem_332 = _RAND_332[255:0];
  _RAND_333 = {8{`RANDOM}};
  mem_333 = _RAND_333[255:0];
  _RAND_334 = {8{`RANDOM}};
  mem_334 = _RAND_334[255:0];
  _RAND_335 = {8{`RANDOM}};
  mem_335 = _RAND_335[255:0];
  _RAND_336 = {8{`RANDOM}};
  mem_336 = _RAND_336[255:0];
  _RAND_337 = {8{`RANDOM}};
  mem_337 = _RAND_337[255:0];
  _RAND_338 = {8{`RANDOM}};
  mem_338 = _RAND_338[255:0];
  _RAND_339 = {8{`RANDOM}};
  mem_339 = _RAND_339[255:0];
  _RAND_340 = {8{`RANDOM}};
  mem_340 = _RAND_340[255:0];
  _RAND_341 = {8{`RANDOM}};
  mem_341 = _RAND_341[255:0];
  _RAND_342 = {8{`RANDOM}};
  mem_342 = _RAND_342[255:0];
  _RAND_343 = {8{`RANDOM}};
  mem_343 = _RAND_343[255:0];
  _RAND_344 = {8{`RANDOM}};
  mem_344 = _RAND_344[255:0];
  _RAND_345 = {8{`RANDOM}};
  mem_345 = _RAND_345[255:0];
  _RAND_346 = {8{`RANDOM}};
  mem_346 = _RAND_346[255:0];
  _RAND_347 = {8{`RANDOM}};
  mem_347 = _RAND_347[255:0];
  _RAND_348 = {8{`RANDOM}};
  mem_348 = _RAND_348[255:0];
  _RAND_349 = {8{`RANDOM}};
  mem_349 = _RAND_349[255:0];
  _RAND_350 = {8{`RANDOM}};
  mem_350 = _RAND_350[255:0];
  _RAND_351 = {8{`RANDOM}};
  mem_351 = _RAND_351[255:0];
  _RAND_352 = {8{`RANDOM}};
  mem_352 = _RAND_352[255:0];
  _RAND_353 = {8{`RANDOM}};
  mem_353 = _RAND_353[255:0];
  _RAND_354 = {8{`RANDOM}};
  mem_354 = _RAND_354[255:0];
  _RAND_355 = {8{`RANDOM}};
  mem_355 = _RAND_355[255:0];
  _RAND_356 = {8{`RANDOM}};
  mem_356 = _RAND_356[255:0];
  _RAND_357 = {8{`RANDOM}};
  mem_357 = _RAND_357[255:0];
  _RAND_358 = {8{`RANDOM}};
  mem_358 = _RAND_358[255:0];
  _RAND_359 = {8{`RANDOM}};
  mem_359 = _RAND_359[255:0];
  _RAND_360 = {8{`RANDOM}};
  mem_360 = _RAND_360[255:0];
  _RAND_361 = {8{`RANDOM}};
  mem_361 = _RAND_361[255:0];
  _RAND_362 = {8{`RANDOM}};
  mem_362 = _RAND_362[255:0];
  _RAND_363 = {8{`RANDOM}};
  mem_363 = _RAND_363[255:0];
  _RAND_364 = {8{`RANDOM}};
  mem_364 = _RAND_364[255:0];
  _RAND_365 = {8{`RANDOM}};
  mem_365 = _RAND_365[255:0];
  _RAND_366 = {8{`RANDOM}};
  mem_366 = _RAND_366[255:0];
  _RAND_367 = {8{`RANDOM}};
  mem_367 = _RAND_367[255:0];
  _RAND_368 = {8{`RANDOM}};
  mem_368 = _RAND_368[255:0];
  _RAND_369 = {8{`RANDOM}};
  mem_369 = _RAND_369[255:0];
  _RAND_370 = {8{`RANDOM}};
  mem_370 = _RAND_370[255:0];
  _RAND_371 = {8{`RANDOM}};
  mem_371 = _RAND_371[255:0];
  _RAND_372 = {8{`RANDOM}};
  mem_372 = _RAND_372[255:0];
  _RAND_373 = {8{`RANDOM}};
  mem_373 = _RAND_373[255:0];
  _RAND_374 = {8{`RANDOM}};
  mem_374 = _RAND_374[255:0];
  _RAND_375 = {8{`RANDOM}};
  mem_375 = _RAND_375[255:0];
  _RAND_376 = {8{`RANDOM}};
  mem_376 = _RAND_376[255:0];
  _RAND_377 = {8{`RANDOM}};
  mem_377 = _RAND_377[255:0];
  _RAND_378 = {8{`RANDOM}};
  mem_378 = _RAND_378[255:0];
  _RAND_379 = {8{`RANDOM}};
  mem_379 = _RAND_379[255:0];
  _RAND_380 = {8{`RANDOM}};
  mem_380 = _RAND_380[255:0];
  _RAND_381 = {8{`RANDOM}};
  mem_381 = _RAND_381[255:0];
  _RAND_382 = {8{`RANDOM}};
  mem_382 = _RAND_382[255:0];
  _RAND_383 = {8{`RANDOM}};
  mem_383 = _RAND_383[255:0];
  _RAND_384 = {8{`RANDOM}};
  mem_384 = _RAND_384[255:0];
  _RAND_385 = {8{`RANDOM}};
  mem_385 = _RAND_385[255:0];
  _RAND_386 = {8{`RANDOM}};
  mem_386 = _RAND_386[255:0];
  _RAND_387 = {8{`RANDOM}};
  mem_387 = _RAND_387[255:0];
  _RAND_388 = {8{`RANDOM}};
  mem_388 = _RAND_388[255:0];
  _RAND_389 = {8{`RANDOM}};
  mem_389 = _RAND_389[255:0];
  _RAND_390 = {8{`RANDOM}};
  mem_390 = _RAND_390[255:0];
  _RAND_391 = {8{`RANDOM}};
  mem_391 = _RAND_391[255:0];
  _RAND_392 = {8{`RANDOM}};
  mem_392 = _RAND_392[255:0];
  _RAND_393 = {8{`RANDOM}};
  mem_393 = _RAND_393[255:0];
  _RAND_394 = {8{`RANDOM}};
  mem_394 = _RAND_394[255:0];
  _RAND_395 = {8{`RANDOM}};
  mem_395 = _RAND_395[255:0];
  _RAND_396 = {8{`RANDOM}};
  mem_396 = _RAND_396[255:0];
  _RAND_397 = {8{`RANDOM}};
  mem_397 = _RAND_397[255:0];
  _RAND_398 = {8{`RANDOM}};
  mem_398 = _RAND_398[255:0];
  _RAND_399 = {8{`RANDOM}};
  mem_399 = _RAND_399[255:0];
  _RAND_400 = {8{`RANDOM}};
  mem_400 = _RAND_400[255:0];
  _RAND_401 = {8{`RANDOM}};
  mem_401 = _RAND_401[255:0];
  _RAND_402 = {8{`RANDOM}};
  mem_402 = _RAND_402[255:0];
  _RAND_403 = {8{`RANDOM}};
  mem_403 = _RAND_403[255:0];
  _RAND_404 = {8{`RANDOM}};
  mem_404 = _RAND_404[255:0];
  _RAND_405 = {8{`RANDOM}};
  mem_405 = _RAND_405[255:0];
  _RAND_406 = {8{`RANDOM}};
  mem_406 = _RAND_406[255:0];
  _RAND_407 = {8{`RANDOM}};
  mem_407 = _RAND_407[255:0];
  _RAND_408 = {8{`RANDOM}};
  mem_408 = _RAND_408[255:0];
  _RAND_409 = {8{`RANDOM}};
  mem_409 = _RAND_409[255:0];
  _RAND_410 = {8{`RANDOM}};
  mem_410 = _RAND_410[255:0];
  _RAND_411 = {8{`RANDOM}};
  mem_411 = _RAND_411[255:0];
  _RAND_412 = {8{`RANDOM}};
  mem_412 = _RAND_412[255:0];
  _RAND_413 = {8{`RANDOM}};
  mem_413 = _RAND_413[255:0];
  _RAND_414 = {8{`RANDOM}};
  mem_414 = _RAND_414[255:0];
  _RAND_415 = {8{`RANDOM}};
  mem_415 = _RAND_415[255:0];
  _RAND_416 = {8{`RANDOM}};
  mem_416 = _RAND_416[255:0];
  _RAND_417 = {8{`RANDOM}};
  mem_417 = _RAND_417[255:0];
  _RAND_418 = {8{`RANDOM}};
  mem_418 = _RAND_418[255:0];
  _RAND_419 = {8{`RANDOM}};
  mem_419 = _RAND_419[255:0];
  _RAND_420 = {8{`RANDOM}};
  mem_420 = _RAND_420[255:0];
  _RAND_421 = {8{`RANDOM}};
  mem_421 = _RAND_421[255:0];
  _RAND_422 = {8{`RANDOM}};
  mem_422 = _RAND_422[255:0];
  _RAND_423 = {8{`RANDOM}};
  mem_423 = _RAND_423[255:0];
  _RAND_424 = {8{`RANDOM}};
  mem_424 = _RAND_424[255:0];
  _RAND_425 = {8{`RANDOM}};
  mem_425 = _RAND_425[255:0];
  _RAND_426 = {8{`RANDOM}};
  mem_426 = _RAND_426[255:0];
  _RAND_427 = {8{`RANDOM}};
  mem_427 = _RAND_427[255:0];
  _RAND_428 = {8{`RANDOM}};
  mem_428 = _RAND_428[255:0];
  _RAND_429 = {8{`RANDOM}};
  mem_429 = _RAND_429[255:0];
  _RAND_430 = {8{`RANDOM}};
  mem_430 = _RAND_430[255:0];
  _RAND_431 = {8{`RANDOM}};
  mem_431 = _RAND_431[255:0];
  _RAND_432 = {8{`RANDOM}};
  mem_432 = _RAND_432[255:0];
  _RAND_433 = {8{`RANDOM}};
  mem_433 = _RAND_433[255:0];
  _RAND_434 = {8{`RANDOM}};
  mem_434 = _RAND_434[255:0];
  _RAND_435 = {8{`RANDOM}};
  mem_435 = _RAND_435[255:0];
  _RAND_436 = {8{`RANDOM}};
  mem_436 = _RAND_436[255:0];
  _RAND_437 = {8{`RANDOM}};
  mem_437 = _RAND_437[255:0];
  _RAND_438 = {8{`RANDOM}};
  mem_438 = _RAND_438[255:0];
  _RAND_439 = {8{`RANDOM}};
  mem_439 = _RAND_439[255:0];
  _RAND_440 = {8{`RANDOM}};
  mem_440 = _RAND_440[255:0];
  _RAND_441 = {8{`RANDOM}};
  mem_441 = _RAND_441[255:0];
  _RAND_442 = {8{`RANDOM}};
  mem_442 = _RAND_442[255:0];
  _RAND_443 = {8{`RANDOM}};
  mem_443 = _RAND_443[255:0];
  _RAND_444 = {8{`RANDOM}};
  mem_444 = _RAND_444[255:0];
  _RAND_445 = {8{`RANDOM}};
  mem_445 = _RAND_445[255:0];
  _RAND_446 = {8{`RANDOM}};
  mem_446 = _RAND_446[255:0];
  _RAND_447 = {8{`RANDOM}};
  mem_447 = _RAND_447[255:0];
  _RAND_448 = {8{`RANDOM}};
  mem_448 = _RAND_448[255:0];
  _RAND_449 = {8{`RANDOM}};
  mem_449 = _RAND_449[255:0];
  _RAND_450 = {8{`RANDOM}};
  mem_450 = _RAND_450[255:0];
  _RAND_451 = {8{`RANDOM}};
  mem_451 = _RAND_451[255:0];
  _RAND_452 = {8{`RANDOM}};
  mem_452 = _RAND_452[255:0];
  _RAND_453 = {8{`RANDOM}};
  mem_453 = _RAND_453[255:0];
  _RAND_454 = {8{`RANDOM}};
  mem_454 = _RAND_454[255:0];
  _RAND_455 = {8{`RANDOM}};
  mem_455 = _RAND_455[255:0];
  _RAND_456 = {8{`RANDOM}};
  mem_456 = _RAND_456[255:0];
  _RAND_457 = {8{`RANDOM}};
  mem_457 = _RAND_457[255:0];
  _RAND_458 = {8{`RANDOM}};
  mem_458 = _RAND_458[255:0];
  _RAND_459 = {8{`RANDOM}};
  mem_459 = _RAND_459[255:0];
  _RAND_460 = {8{`RANDOM}};
  mem_460 = _RAND_460[255:0];
  _RAND_461 = {8{`RANDOM}};
  mem_461 = _RAND_461[255:0];
  _RAND_462 = {8{`RANDOM}};
  mem_462 = _RAND_462[255:0];
  _RAND_463 = {8{`RANDOM}};
  mem_463 = _RAND_463[255:0];
  _RAND_464 = {8{`RANDOM}};
  mem_464 = _RAND_464[255:0];
  _RAND_465 = {8{`RANDOM}};
  mem_465 = _RAND_465[255:0];
  _RAND_466 = {8{`RANDOM}};
  mem_466 = _RAND_466[255:0];
  _RAND_467 = {8{`RANDOM}};
  mem_467 = _RAND_467[255:0];
  _RAND_468 = {8{`RANDOM}};
  mem_468 = _RAND_468[255:0];
  _RAND_469 = {8{`RANDOM}};
  mem_469 = _RAND_469[255:0];
  _RAND_470 = {8{`RANDOM}};
  mem_470 = _RAND_470[255:0];
  _RAND_471 = {8{`RANDOM}};
  mem_471 = _RAND_471[255:0];
  _RAND_472 = {8{`RANDOM}};
  mem_472 = _RAND_472[255:0];
  _RAND_473 = {8{`RANDOM}};
  mem_473 = _RAND_473[255:0];
  _RAND_474 = {8{`RANDOM}};
  mem_474 = _RAND_474[255:0];
  _RAND_475 = {8{`RANDOM}};
  mem_475 = _RAND_475[255:0];
  _RAND_476 = {8{`RANDOM}};
  mem_476 = _RAND_476[255:0];
  _RAND_477 = {8{`RANDOM}};
  mem_477 = _RAND_477[255:0];
  _RAND_478 = {8{`RANDOM}};
  mem_478 = _RAND_478[255:0];
  _RAND_479 = {8{`RANDOM}};
  mem_479 = _RAND_479[255:0];
  _RAND_480 = {8{`RANDOM}};
  mem_480 = _RAND_480[255:0];
  _RAND_481 = {8{`RANDOM}};
  mem_481 = _RAND_481[255:0];
  _RAND_482 = {8{`RANDOM}};
  mem_482 = _RAND_482[255:0];
  _RAND_483 = {8{`RANDOM}};
  mem_483 = _RAND_483[255:0];
  _RAND_484 = {8{`RANDOM}};
  mem_484 = _RAND_484[255:0];
  _RAND_485 = {8{`RANDOM}};
  mem_485 = _RAND_485[255:0];
  _RAND_486 = {8{`RANDOM}};
  mem_486 = _RAND_486[255:0];
  _RAND_487 = {8{`RANDOM}};
  mem_487 = _RAND_487[255:0];
  _RAND_488 = {8{`RANDOM}};
  mem_488 = _RAND_488[255:0];
  _RAND_489 = {8{`RANDOM}};
  mem_489 = _RAND_489[255:0];
  _RAND_490 = {8{`RANDOM}};
  mem_490 = _RAND_490[255:0];
  _RAND_491 = {8{`RANDOM}};
  mem_491 = _RAND_491[255:0];
  _RAND_492 = {8{`RANDOM}};
  mem_492 = _RAND_492[255:0];
  _RAND_493 = {8{`RANDOM}};
  mem_493 = _RAND_493[255:0];
  _RAND_494 = {8{`RANDOM}};
  mem_494 = _RAND_494[255:0];
  _RAND_495 = {8{`RANDOM}};
  mem_495 = _RAND_495[255:0];
  _RAND_496 = {8{`RANDOM}};
  mem_496 = _RAND_496[255:0];
  _RAND_497 = {8{`RANDOM}};
  mem_497 = _RAND_497[255:0];
  _RAND_498 = {8{`RANDOM}};
  mem_498 = _RAND_498[255:0];
  _RAND_499 = {8{`RANDOM}};
  mem_499 = _RAND_499[255:0];
  _RAND_500 = {8{`RANDOM}};
  mem_500 = _RAND_500[255:0];
  _RAND_501 = {8{`RANDOM}};
  mem_501 = _RAND_501[255:0];
  _RAND_502 = {8{`RANDOM}};
  mem_502 = _RAND_502[255:0];
  _RAND_503 = {8{`RANDOM}};
  mem_503 = _RAND_503[255:0];
  _RAND_504 = {8{`RANDOM}};
  mem_504 = _RAND_504[255:0];
  _RAND_505 = {8{`RANDOM}};
  mem_505 = _RAND_505[255:0];
  _RAND_506 = {8{`RANDOM}};
  mem_506 = _RAND_506[255:0];
  _RAND_507 = {8{`RANDOM}};
  mem_507 = _RAND_507[255:0];
  _RAND_508 = {8{`RANDOM}};
  mem_508 = _RAND_508[255:0];
  _RAND_509 = {8{`RANDOM}};
  mem_509 = _RAND_509[255:0];
  _RAND_510 = {8{`RANDOM}};
  mem_510 = _RAND_510[255:0];
  _RAND_511 = {8{`RANDOM}};
  mem_511 = _RAND_511[255:0];
  _RAND_512 = {8{`RANDOM}};
  mem_512 = _RAND_512[255:0];
  _RAND_513 = {8{`RANDOM}};
  mem_513 = _RAND_513[255:0];
  _RAND_514 = {8{`RANDOM}};
  mem_514 = _RAND_514[255:0];
  _RAND_515 = {8{`RANDOM}};
  mem_515 = _RAND_515[255:0];
  _RAND_516 = {8{`RANDOM}};
  mem_516 = _RAND_516[255:0];
  _RAND_517 = {8{`RANDOM}};
  mem_517 = _RAND_517[255:0];
  _RAND_518 = {8{`RANDOM}};
  mem_518 = _RAND_518[255:0];
  _RAND_519 = {8{`RANDOM}};
  mem_519 = _RAND_519[255:0];
  _RAND_520 = {8{`RANDOM}};
  mem_520 = _RAND_520[255:0];
  _RAND_521 = {8{`RANDOM}};
  mem_521 = _RAND_521[255:0];
  _RAND_522 = {8{`RANDOM}};
  mem_522 = _RAND_522[255:0];
  _RAND_523 = {8{`RANDOM}};
  mem_523 = _RAND_523[255:0];
  _RAND_524 = {8{`RANDOM}};
  mem_524 = _RAND_524[255:0];
  _RAND_525 = {8{`RANDOM}};
  mem_525 = _RAND_525[255:0];
  _RAND_526 = {8{`RANDOM}};
  mem_526 = _RAND_526[255:0];
  _RAND_527 = {8{`RANDOM}};
  mem_527 = _RAND_527[255:0];
  _RAND_528 = {8{`RANDOM}};
  mem_528 = _RAND_528[255:0];
  _RAND_529 = {8{`RANDOM}};
  mem_529 = _RAND_529[255:0];
  _RAND_530 = {8{`RANDOM}};
  mem_530 = _RAND_530[255:0];
  _RAND_531 = {8{`RANDOM}};
  mem_531 = _RAND_531[255:0];
  _RAND_532 = {8{`RANDOM}};
  mem_532 = _RAND_532[255:0];
  _RAND_533 = {8{`RANDOM}};
  mem_533 = _RAND_533[255:0];
  _RAND_534 = {8{`RANDOM}};
  mem_534 = _RAND_534[255:0];
  _RAND_535 = {8{`RANDOM}};
  mem_535 = _RAND_535[255:0];
  _RAND_536 = {8{`RANDOM}};
  mem_536 = _RAND_536[255:0];
  _RAND_537 = {8{`RANDOM}};
  mem_537 = _RAND_537[255:0];
  _RAND_538 = {8{`RANDOM}};
  mem_538 = _RAND_538[255:0];
  _RAND_539 = {8{`RANDOM}};
  mem_539 = _RAND_539[255:0];
  _RAND_540 = {8{`RANDOM}};
  mem_540 = _RAND_540[255:0];
  _RAND_541 = {8{`RANDOM}};
  mem_541 = _RAND_541[255:0];
  _RAND_542 = {8{`RANDOM}};
  mem_542 = _RAND_542[255:0];
  _RAND_543 = {8{`RANDOM}};
  mem_543 = _RAND_543[255:0];
  _RAND_544 = {8{`RANDOM}};
  mem_544 = _RAND_544[255:0];
  _RAND_545 = {8{`RANDOM}};
  mem_545 = _RAND_545[255:0];
  _RAND_546 = {8{`RANDOM}};
  mem_546 = _RAND_546[255:0];
  _RAND_547 = {8{`RANDOM}};
  mem_547 = _RAND_547[255:0];
  _RAND_548 = {8{`RANDOM}};
  mem_548 = _RAND_548[255:0];
  _RAND_549 = {8{`RANDOM}};
  mem_549 = _RAND_549[255:0];
  _RAND_550 = {8{`RANDOM}};
  mem_550 = _RAND_550[255:0];
  _RAND_551 = {8{`RANDOM}};
  mem_551 = _RAND_551[255:0];
  _RAND_552 = {8{`RANDOM}};
  mem_552 = _RAND_552[255:0];
  _RAND_553 = {8{`RANDOM}};
  mem_553 = _RAND_553[255:0];
  _RAND_554 = {8{`RANDOM}};
  mem_554 = _RAND_554[255:0];
  _RAND_555 = {8{`RANDOM}};
  mem_555 = _RAND_555[255:0];
  _RAND_556 = {8{`RANDOM}};
  mem_556 = _RAND_556[255:0];
  _RAND_557 = {8{`RANDOM}};
  mem_557 = _RAND_557[255:0];
  _RAND_558 = {8{`RANDOM}};
  mem_558 = _RAND_558[255:0];
  _RAND_559 = {8{`RANDOM}};
  mem_559 = _RAND_559[255:0];
  _RAND_560 = {8{`RANDOM}};
  mem_560 = _RAND_560[255:0];
  _RAND_561 = {8{`RANDOM}};
  mem_561 = _RAND_561[255:0];
  _RAND_562 = {8{`RANDOM}};
  mem_562 = _RAND_562[255:0];
  _RAND_563 = {8{`RANDOM}};
  mem_563 = _RAND_563[255:0];
  _RAND_564 = {8{`RANDOM}};
  mem_564 = _RAND_564[255:0];
  _RAND_565 = {8{`RANDOM}};
  mem_565 = _RAND_565[255:0];
  _RAND_566 = {8{`RANDOM}};
  mem_566 = _RAND_566[255:0];
  _RAND_567 = {8{`RANDOM}};
  mem_567 = _RAND_567[255:0];
  _RAND_568 = {8{`RANDOM}};
  mem_568 = _RAND_568[255:0];
  _RAND_569 = {8{`RANDOM}};
  mem_569 = _RAND_569[255:0];
  _RAND_570 = {8{`RANDOM}};
  mem_570 = _RAND_570[255:0];
  _RAND_571 = {8{`RANDOM}};
  mem_571 = _RAND_571[255:0];
  _RAND_572 = {8{`RANDOM}};
  mem_572 = _RAND_572[255:0];
  _RAND_573 = {8{`RANDOM}};
  mem_573 = _RAND_573[255:0];
  _RAND_574 = {8{`RANDOM}};
  mem_574 = _RAND_574[255:0];
  _RAND_575 = {8{`RANDOM}};
  mem_575 = _RAND_575[255:0];
  _RAND_576 = {8{`RANDOM}};
  mem_576 = _RAND_576[255:0];
  _RAND_577 = {8{`RANDOM}};
  mem_577 = _RAND_577[255:0];
  _RAND_578 = {8{`RANDOM}};
  mem_578 = _RAND_578[255:0];
  _RAND_579 = {8{`RANDOM}};
  mem_579 = _RAND_579[255:0];
  _RAND_580 = {8{`RANDOM}};
  mem_580 = _RAND_580[255:0];
  _RAND_581 = {8{`RANDOM}};
  mem_581 = _RAND_581[255:0];
  _RAND_582 = {8{`RANDOM}};
  mem_582 = _RAND_582[255:0];
  _RAND_583 = {8{`RANDOM}};
  mem_583 = _RAND_583[255:0];
  _RAND_584 = {8{`RANDOM}};
  mem_584 = _RAND_584[255:0];
  _RAND_585 = {8{`RANDOM}};
  mem_585 = _RAND_585[255:0];
  _RAND_586 = {8{`RANDOM}};
  mem_586 = _RAND_586[255:0];
  _RAND_587 = {8{`RANDOM}};
  mem_587 = _RAND_587[255:0];
  _RAND_588 = {8{`RANDOM}};
  mem_588 = _RAND_588[255:0];
  _RAND_589 = {8{`RANDOM}};
  mem_589 = _RAND_589[255:0];
  _RAND_590 = {8{`RANDOM}};
  mem_590 = _RAND_590[255:0];
  _RAND_591 = {8{`RANDOM}};
  mem_591 = _RAND_591[255:0];
  _RAND_592 = {8{`RANDOM}};
  mem_592 = _RAND_592[255:0];
  _RAND_593 = {8{`RANDOM}};
  mem_593 = _RAND_593[255:0];
  _RAND_594 = {8{`RANDOM}};
  mem_594 = _RAND_594[255:0];
  _RAND_595 = {8{`RANDOM}};
  mem_595 = _RAND_595[255:0];
  _RAND_596 = {8{`RANDOM}};
  mem_596 = _RAND_596[255:0];
  _RAND_597 = {8{`RANDOM}};
  mem_597 = _RAND_597[255:0];
  _RAND_598 = {8{`RANDOM}};
  mem_598 = _RAND_598[255:0];
  _RAND_599 = {8{`RANDOM}};
  mem_599 = _RAND_599[255:0];
  _RAND_600 = {8{`RANDOM}};
  mem_600 = _RAND_600[255:0];
  _RAND_601 = {8{`RANDOM}};
  mem_601 = _RAND_601[255:0];
  _RAND_602 = {8{`RANDOM}};
  mem_602 = _RAND_602[255:0];
  _RAND_603 = {8{`RANDOM}};
  mem_603 = _RAND_603[255:0];
  _RAND_604 = {8{`RANDOM}};
  mem_604 = _RAND_604[255:0];
  _RAND_605 = {8{`RANDOM}};
  mem_605 = _RAND_605[255:0];
  _RAND_606 = {8{`RANDOM}};
  mem_606 = _RAND_606[255:0];
  _RAND_607 = {8{`RANDOM}};
  mem_607 = _RAND_607[255:0];
  _RAND_608 = {8{`RANDOM}};
  mem_608 = _RAND_608[255:0];
  _RAND_609 = {8{`RANDOM}};
  mem_609 = _RAND_609[255:0];
  _RAND_610 = {8{`RANDOM}};
  mem_610 = _RAND_610[255:0];
  _RAND_611 = {8{`RANDOM}};
  mem_611 = _RAND_611[255:0];
  _RAND_612 = {8{`RANDOM}};
  mem_612 = _RAND_612[255:0];
  _RAND_613 = {8{`RANDOM}};
  mem_613 = _RAND_613[255:0];
  _RAND_614 = {8{`RANDOM}};
  mem_614 = _RAND_614[255:0];
  _RAND_615 = {8{`RANDOM}};
  mem_615 = _RAND_615[255:0];
  _RAND_616 = {8{`RANDOM}};
  mem_616 = _RAND_616[255:0];
  _RAND_617 = {8{`RANDOM}};
  mem_617 = _RAND_617[255:0];
  _RAND_618 = {8{`RANDOM}};
  mem_618 = _RAND_618[255:0];
  _RAND_619 = {8{`RANDOM}};
  mem_619 = _RAND_619[255:0];
  _RAND_620 = {8{`RANDOM}};
  mem_620 = _RAND_620[255:0];
  _RAND_621 = {8{`RANDOM}};
  mem_621 = _RAND_621[255:0];
  _RAND_622 = {8{`RANDOM}};
  mem_622 = _RAND_622[255:0];
  _RAND_623 = {8{`RANDOM}};
  mem_623 = _RAND_623[255:0];
  _RAND_624 = {8{`RANDOM}};
  mem_624 = _RAND_624[255:0];
  _RAND_625 = {8{`RANDOM}};
  mem_625 = _RAND_625[255:0];
  _RAND_626 = {8{`RANDOM}};
  mem_626 = _RAND_626[255:0];
  _RAND_627 = {8{`RANDOM}};
  mem_627 = _RAND_627[255:0];
  _RAND_628 = {8{`RANDOM}};
  mem_628 = _RAND_628[255:0];
  _RAND_629 = {8{`RANDOM}};
  mem_629 = _RAND_629[255:0];
  _RAND_630 = {8{`RANDOM}};
  mem_630 = _RAND_630[255:0];
  _RAND_631 = {8{`RANDOM}};
  mem_631 = _RAND_631[255:0];
  _RAND_632 = {8{`RANDOM}};
  mem_632 = _RAND_632[255:0];
  _RAND_633 = {8{`RANDOM}};
  mem_633 = _RAND_633[255:0];
  _RAND_634 = {8{`RANDOM}};
  mem_634 = _RAND_634[255:0];
  _RAND_635 = {8{`RANDOM}};
  mem_635 = _RAND_635[255:0];
  _RAND_636 = {8{`RANDOM}};
  mem_636 = _RAND_636[255:0];
  _RAND_637 = {8{`RANDOM}};
  mem_637 = _RAND_637[255:0];
  _RAND_638 = {8{`RANDOM}};
  mem_638 = _RAND_638[255:0];
  _RAND_639 = {8{`RANDOM}};
  mem_639 = _RAND_639[255:0];
  _RAND_640 = {8{`RANDOM}};
  mem_640 = _RAND_640[255:0];
  _RAND_641 = {8{`RANDOM}};
  mem_641 = _RAND_641[255:0];
  _RAND_642 = {8{`RANDOM}};
  mem_642 = _RAND_642[255:0];
  _RAND_643 = {8{`RANDOM}};
  mem_643 = _RAND_643[255:0];
  _RAND_644 = {8{`RANDOM}};
  mem_644 = _RAND_644[255:0];
  _RAND_645 = {8{`RANDOM}};
  mem_645 = _RAND_645[255:0];
  _RAND_646 = {8{`RANDOM}};
  mem_646 = _RAND_646[255:0];
  _RAND_647 = {8{`RANDOM}};
  mem_647 = _RAND_647[255:0];
  _RAND_648 = {8{`RANDOM}};
  mem_648 = _RAND_648[255:0];
  _RAND_649 = {8{`RANDOM}};
  mem_649 = _RAND_649[255:0];
  _RAND_650 = {8{`RANDOM}};
  mem_650 = _RAND_650[255:0];
  _RAND_651 = {8{`RANDOM}};
  mem_651 = _RAND_651[255:0];
  _RAND_652 = {8{`RANDOM}};
  mem_652 = _RAND_652[255:0];
  _RAND_653 = {8{`RANDOM}};
  mem_653 = _RAND_653[255:0];
  _RAND_654 = {8{`RANDOM}};
  mem_654 = _RAND_654[255:0];
  _RAND_655 = {8{`RANDOM}};
  mem_655 = _RAND_655[255:0];
  _RAND_656 = {8{`RANDOM}};
  mem_656 = _RAND_656[255:0];
  _RAND_657 = {8{`RANDOM}};
  mem_657 = _RAND_657[255:0];
  _RAND_658 = {8{`RANDOM}};
  mem_658 = _RAND_658[255:0];
  _RAND_659 = {8{`RANDOM}};
  mem_659 = _RAND_659[255:0];
  _RAND_660 = {8{`RANDOM}};
  mem_660 = _RAND_660[255:0];
  _RAND_661 = {8{`RANDOM}};
  mem_661 = _RAND_661[255:0];
  _RAND_662 = {8{`RANDOM}};
  mem_662 = _RAND_662[255:0];
  _RAND_663 = {8{`RANDOM}};
  mem_663 = _RAND_663[255:0];
  _RAND_664 = {8{`RANDOM}};
  mem_664 = _RAND_664[255:0];
  _RAND_665 = {8{`RANDOM}};
  mem_665 = _RAND_665[255:0];
  _RAND_666 = {8{`RANDOM}};
  mem_666 = _RAND_666[255:0];
  _RAND_667 = {8{`RANDOM}};
  mem_667 = _RAND_667[255:0];
  _RAND_668 = {8{`RANDOM}};
  mem_668 = _RAND_668[255:0];
  _RAND_669 = {8{`RANDOM}};
  mem_669 = _RAND_669[255:0];
  _RAND_670 = {8{`RANDOM}};
  mem_670 = _RAND_670[255:0];
  _RAND_671 = {8{`RANDOM}};
  mem_671 = _RAND_671[255:0];
  _RAND_672 = {8{`RANDOM}};
  mem_672 = _RAND_672[255:0];
  _RAND_673 = {8{`RANDOM}};
  mem_673 = _RAND_673[255:0];
  _RAND_674 = {8{`RANDOM}};
  mem_674 = _RAND_674[255:0];
  _RAND_675 = {8{`RANDOM}};
  mem_675 = _RAND_675[255:0];
  _RAND_676 = {8{`RANDOM}};
  mem_676 = _RAND_676[255:0];
  _RAND_677 = {8{`RANDOM}};
  mem_677 = _RAND_677[255:0];
  _RAND_678 = {8{`RANDOM}};
  mem_678 = _RAND_678[255:0];
  _RAND_679 = {8{`RANDOM}};
  mem_679 = _RAND_679[255:0];
  _RAND_680 = {8{`RANDOM}};
  mem_680 = _RAND_680[255:0];
  _RAND_681 = {8{`RANDOM}};
  mem_681 = _RAND_681[255:0];
  _RAND_682 = {8{`RANDOM}};
  mem_682 = _RAND_682[255:0];
  _RAND_683 = {8{`RANDOM}};
  mem_683 = _RAND_683[255:0];
  _RAND_684 = {8{`RANDOM}};
  mem_684 = _RAND_684[255:0];
  _RAND_685 = {8{`RANDOM}};
  mem_685 = _RAND_685[255:0];
  _RAND_686 = {8{`RANDOM}};
  mem_686 = _RAND_686[255:0];
  _RAND_687 = {8{`RANDOM}};
  mem_687 = _RAND_687[255:0];
  _RAND_688 = {8{`RANDOM}};
  mem_688 = _RAND_688[255:0];
  _RAND_689 = {8{`RANDOM}};
  mem_689 = _RAND_689[255:0];
  _RAND_690 = {8{`RANDOM}};
  mem_690 = _RAND_690[255:0];
  _RAND_691 = {8{`RANDOM}};
  mem_691 = _RAND_691[255:0];
  _RAND_692 = {8{`RANDOM}};
  mem_692 = _RAND_692[255:0];
  _RAND_693 = {8{`RANDOM}};
  mem_693 = _RAND_693[255:0];
  _RAND_694 = {8{`RANDOM}};
  mem_694 = _RAND_694[255:0];
  _RAND_695 = {8{`RANDOM}};
  mem_695 = _RAND_695[255:0];
  _RAND_696 = {8{`RANDOM}};
  mem_696 = _RAND_696[255:0];
  _RAND_697 = {8{`RANDOM}};
  mem_697 = _RAND_697[255:0];
  _RAND_698 = {8{`RANDOM}};
  mem_698 = _RAND_698[255:0];
  _RAND_699 = {8{`RANDOM}};
  mem_699 = _RAND_699[255:0];
  _RAND_700 = {8{`RANDOM}};
  mem_700 = _RAND_700[255:0];
  _RAND_701 = {8{`RANDOM}};
  mem_701 = _RAND_701[255:0];
  _RAND_702 = {8{`RANDOM}};
  mem_702 = _RAND_702[255:0];
  _RAND_703 = {8{`RANDOM}};
  mem_703 = _RAND_703[255:0];
  _RAND_704 = {8{`RANDOM}};
  mem_704 = _RAND_704[255:0];
  _RAND_705 = {8{`RANDOM}};
  mem_705 = _RAND_705[255:0];
  _RAND_706 = {8{`RANDOM}};
  mem_706 = _RAND_706[255:0];
  _RAND_707 = {8{`RANDOM}};
  mem_707 = _RAND_707[255:0];
  _RAND_708 = {8{`RANDOM}};
  mem_708 = _RAND_708[255:0];
  _RAND_709 = {8{`RANDOM}};
  mem_709 = _RAND_709[255:0];
  _RAND_710 = {8{`RANDOM}};
  mem_710 = _RAND_710[255:0];
  _RAND_711 = {8{`RANDOM}};
  mem_711 = _RAND_711[255:0];
  _RAND_712 = {8{`RANDOM}};
  mem_712 = _RAND_712[255:0];
  _RAND_713 = {8{`RANDOM}};
  mem_713 = _RAND_713[255:0];
  _RAND_714 = {8{`RANDOM}};
  mem_714 = _RAND_714[255:0];
  _RAND_715 = {8{`RANDOM}};
  mem_715 = _RAND_715[255:0];
  _RAND_716 = {8{`RANDOM}};
  mem_716 = _RAND_716[255:0];
  _RAND_717 = {8{`RANDOM}};
  mem_717 = _RAND_717[255:0];
  _RAND_718 = {8{`RANDOM}};
  mem_718 = _RAND_718[255:0];
  _RAND_719 = {8{`RANDOM}};
  mem_719 = _RAND_719[255:0];
  _RAND_720 = {8{`RANDOM}};
  mem_720 = _RAND_720[255:0];
  _RAND_721 = {8{`RANDOM}};
  mem_721 = _RAND_721[255:0];
  _RAND_722 = {8{`RANDOM}};
  mem_722 = _RAND_722[255:0];
  _RAND_723 = {8{`RANDOM}};
  mem_723 = _RAND_723[255:0];
  _RAND_724 = {8{`RANDOM}};
  mem_724 = _RAND_724[255:0];
  _RAND_725 = {8{`RANDOM}};
  mem_725 = _RAND_725[255:0];
  _RAND_726 = {8{`RANDOM}};
  mem_726 = _RAND_726[255:0];
  _RAND_727 = {8{`RANDOM}};
  mem_727 = _RAND_727[255:0];
  _RAND_728 = {8{`RANDOM}};
  mem_728 = _RAND_728[255:0];
  _RAND_729 = {8{`RANDOM}};
  mem_729 = _RAND_729[255:0];
  _RAND_730 = {8{`RANDOM}};
  mem_730 = _RAND_730[255:0];
  _RAND_731 = {8{`RANDOM}};
  mem_731 = _RAND_731[255:0];
  _RAND_732 = {8{`RANDOM}};
  mem_732 = _RAND_732[255:0];
  _RAND_733 = {8{`RANDOM}};
  mem_733 = _RAND_733[255:0];
  _RAND_734 = {8{`RANDOM}};
  mem_734 = _RAND_734[255:0];
  _RAND_735 = {8{`RANDOM}};
  mem_735 = _RAND_735[255:0];
  _RAND_736 = {8{`RANDOM}};
  mem_736 = _RAND_736[255:0];
  _RAND_737 = {8{`RANDOM}};
  mem_737 = _RAND_737[255:0];
  _RAND_738 = {8{`RANDOM}};
  mem_738 = _RAND_738[255:0];
  _RAND_739 = {8{`RANDOM}};
  mem_739 = _RAND_739[255:0];
  _RAND_740 = {8{`RANDOM}};
  mem_740 = _RAND_740[255:0];
  _RAND_741 = {8{`RANDOM}};
  mem_741 = _RAND_741[255:0];
  _RAND_742 = {8{`RANDOM}};
  mem_742 = _RAND_742[255:0];
  _RAND_743 = {8{`RANDOM}};
  mem_743 = _RAND_743[255:0];
  _RAND_744 = {8{`RANDOM}};
  mem_744 = _RAND_744[255:0];
  _RAND_745 = {8{`RANDOM}};
  mem_745 = _RAND_745[255:0];
  _RAND_746 = {8{`RANDOM}};
  mem_746 = _RAND_746[255:0];
  _RAND_747 = {8{`RANDOM}};
  mem_747 = _RAND_747[255:0];
  _RAND_748 = {8{`RANDOM}};
  mem_748 = _RAND_748[255:0];
  _RAND_749 = {8{`RANDOM}};
  mem_749 = _RAND_749[255:0];
  _RAND_750 = {8{`RANDOM}};
  mem_750 = _RAND_750[255:0];
  _RAND_751 = {8{`RANDOM}};
  mem_751 = _RAND_751[255:0];
  _RAND_752 = {8{`RANDOM}};
  mem_752 = _RAND_752[255:0];
  _RAND_753 = {8{`RANDOM}};
  mem_753 = _RAND_753[255:0];
  _RAND_754 = {8{`RANDOM}};
  mem_754 = _RAND_754[255:0];
  _RAND_755 = {8{`RANDOM}};
  mem_755 = _RAND_755[255:0];
  _RAND_756 = {8{`RANDOM}};
  mem_756 = _RAND_756[255:0];
  _RAND_757 = {8{`RANDOM}};
  mem_757 = _RAND_757[255:0];
  _RAND_758 = {8{`RANDOM}};
  mem_758 = _RAND_758[255:0];
  _RAND_759 = {8{`RANDOM}};
  mem_759 = _RAND_759[255:0];
  _RAND_760 = {8{`RANDOM}};
  mem_760 = _RAND_760[255:0];
  _RAND_761 = {8{`RANDOM}};
  mem_761 = _RAND_761[255:0];
  _RAND_762 = {8{`RANDOM}};
  mem_762 = _RAND_762[255:0];
  _RAND_763 = {8{`RANDOM}};
  mem_763 = _RAND_763[255:0];
  _RAND_764 = {8{`RANDOM}};
  mem_764 = _RAND_764[255:0];
  _RAND_765 = {8{`RANDOM}};
  mem_765 = _RAND_765[255:0];
  _RAND_766 = {8{`RANDOM}};
  mem_766 = _RAND_766[255:0];
  _RAND_767 = {8{`RANDOM}};
  mem_767 = _RAND_767[255:0];
  _RAND_768 = {8{`RANDOM}};
  mem_768 = _RAND_768[255:0];
  _RAND_769 = {8{`RANDOM}};
  mem_769 = _RAND_769[255:0];
  _RAND_770 = {8{`RANDOM}};
  mem_770 = _RAND_770[255:0];
  _RAND_771 = {8{`RANDOM}};
  mem_771 = _RAND_771[255:0];
  _RAND_772 = {8{`RANDOM}};
  mem_772 = _RAND_772[255:0];
  _RAND_773 = {8{`RANDOM}};
  mem_773 = _RAND_773[255:0];
  _RAND_774 = {8{`RANDOM}};
  mem_774 = _RAND_774[255:0];
  _RAND_775 = {8{`RANDOM}};
  mem_775 = _RAND_775[255:0];
  _RAND_776 = {8{`RANDOM}};
  mem_776 = _RAND_776[255:0];
  _RAND_777 = {8{`RANDOM}};
  mem_777 = _RAND_777[255:0];
  _RAND_778 = {8{`RANDOM}};
  mem_778 = _RAND_778[255:0];
  _RAND_779 = {8{`RANDOM}};
  mem_779 = _RAND_779[255:0];
  _RAND_780 = {8{`RANDOM}};
  mem_780 = _RAND_780[255:0];
  _RAND_781 = {8{`RANDOM}};
  mem_781 = _RAND_781[255:0];
  _RAND_782 = {8{`RANDOM}};
  mem_782 = _RAND_782[255:0];
  _RAND_783 = {8{`RANDOM}};
  mem_783 = _RAND_783[255:0];
  _RAND_784 = {8{`RANDOM}};
  mem_784 = _RAND_784[255:0];
  _RAND_785 = {8{`RANDOM}};
  mem_785 = _RAND_785[255:0];
  _RAND_786 = {8{`RANDOM}};
  mem_786 = _RAND_786[255:0];
  _RAND_787 = {8{`RANDOM}};
  mem_787 = _RAND_787[255:0];
  _RAND_788 = {8{`RANDOM}};
  mem_788 = _RAND_788[255:0];
  _RAND_789 = {8{`RANDOM}};
  mem_789 = _RAND_789[255:0];
  _RAND_790 = {8{`RANDOM}};
  mem_790 = _RAND_790[255:0];
  _RAND_791 = {8{`RANDOM}};
  mem_791 = _RAND_791[255:0];
  _RAND_792 = {8{`RANDOM}};
  mem_792 = _RAND_792[255:0];
  _RAND_793 = {8{`RANDOM}};
  mem_793 = _RAND_793[255:0];
  _RAND_794 = {8{`RANDOM}};
  mem_794 = _RAND_794[255:0];
  _RAND_795 = {8{`RANDOM}};
  mem_795 = _RAND_795[255:0];
  _RAND_796 = {8{`RANDOM}};
  mem_796 = _RAND_796[255:0];
  _RAND_797 = {8{`RANDOM}};
  mem_797 = _RAND_797[255:0];
  _RAND_798 = {8{`RANDOM}};
  mem_798 = _RAND_798[255:0];
  _RAND_799 = {8{`RANDOM}};
  mem_799 = _RAND_799[255:0];
  _RAND_800 = {8{`RANDOM}};
  mem_800 = _RAND_800[255:0];
  _RAND_801 = {8{`RANDOM}};
  mem_801 = _RAND_801[255:0];
  _RAND_802 = {8{`RANDOM}};
  mem_802 = _RAND_802[255:0];
  _RAND_803 = {8{`RANDOM}};
  mem_803 = _RAND_803[255:0];
  _RAND_804 = {8{`RANDOM}};
  mem_804 = _RAND_804[255:0];
  _RAND_805 = {8{`RANDOM}};
  mem_805 = _RAND_805[255:0];
  _RAND_806 = {8{`RANDOM}};
  mem_806 = _RAND_806[255:0];
  _RAND_807 = {8{`RANDOM}};
  mem_807 = _RAND_807[255:0];
  _RAND_808 = {8{`RANDOM}};
  mem_808 = _RAND_808[255:0];
  _RAND_809 = {8{`RANDOM}};
  mem_809 = _RAND_809[255:0];
  _RAND_810 = {8{`RANDOM}};
  mem_810 = _RAND_810[255:0];
  _RAND_811 = {8{`RANDOM}};
  mem_811 = _RAND_811[255:0];
  _RAND_812 = {8{`RANDOM}};
  mem_812 = _RAND_812[255:0];
  _RAND_813 = {8{`RANDOM}};
  mem_813 = _RAND_813[255:0];
  _RAND_814 = {8{`RANDOM}};
  mem_814 = _RAND_814[255:0];
  _RAND_815 = {8{`RANDOM}};
  mem_815 = _RAND_815[255:0];
  _RAND_816 = {8{`RANDOM}};
  mem_816 = _RAND_816[255:0];
  _RAND_817 = {8{`RANDOM}};
  mem_817 = _RAND_817[255:0];
  _RAND_818 = {8{`RANDOM}};
  mem_818 = _RAND_818[255:0];
  _RAND_819 = {8{`RANDOM}};
  mem_819 = _RAND_819[255:0];
  _RAND_820 = {8{`RANDOM}};
  mem_820 = _RAND_820[255:0];
  _RAND_821 = {8{`RANDOM}};
  mem_821 = _RAND_821[255:0];
  _RAND_822 = {8{`RANDOM}};
  mem_822 = _RAND_822[255:0];
  _RAND_823 = {8{`RANDOM}};
  mem_823 = _RAND_823[255:0];
  _RAND_824 = {8{`RANDOM}};
  mem_824 = _RAND_824[255:0];
  _RAND_825 = {8{`RANDOM}};
  mem_825 = _RAND_825[255:0];
  _RAND_826 = {8{`RANDOM}};
  mem_826 = _RAND_826[255:0];
  _RAND_827 = {8{`RANDOM}};
  mem_827 = _RAND_827[255:0];
  _RAND_828 = {8{`RANDOM}};
  mem_828 = _RAND_828[255:0];
  _RAND_829 = {8{`RANDOM}};
  mem_829 = _RAND_829[255:0];
  _RAND_830 = {8{`RANDOM}};
  mem_830 = _RAND_830[255:0];
  _RAND_831 = {8{`RANDOM}};
  mem_831 = _RAND_831[255:0];
  _RAND_832 = {8{`RANDOM}};
  mem_832 = _RAND_832[255:0];
  _RAND_833 = {8{`RANDOM}};
  mem_833 = _RAND_833[255:0];
  _RAND_834 = {8{`RANDOM}};
  mem_834 = _RAND_834[255:0];
  _RAND_835 = {8{`RANDOM}};
  mem_835 = _RAND_835[255:0];
  _RAND_836 = {8{`RANDOM}};
  mem_836 = _RAND_836[255:0];
  _RAND_837 = {8{`RANDOM}};
  mem_837 = _RAND_837[255:0];
  _RAND_838 = {8{`RANDOM}};
  mem_838 = _RAND_838[255:0];
  _RAND_839 = {8{`RANDOM}};
  mem_839 = _RAND_839[255:0];
  _RAND_840 = {8{`RANDOM}};
  mem_840 = _RAND_840[255:0];
  _RAND_841 = {8{`RANDOM}};
  mem_841 = _RAND_841[255:0];
  _RAND_842 = {8{`RANDOM}};
  mem_842 = _RAND_842[255:0];
  _RAND_843 = {8{`RANDOM}};
  mem_843 = _RAND_843[255:0];
  _RAND_844 = {8{`RANDOM}};
  mem_844 = _RAND_844[255:0];
  _RAND_845 = {8{`RANDOM}};
  mem_845 = _RAND_845[255:0];
  _RAND_846 = {8{`RANDOM}};
  mem_846 = _RAND_846[255:0];
  _RAND_847 = {8{`RANDOM}};
  mem_847 = _RAND_847[255:0];
  _RAND_848 = {8{`RANDOM}};
  mem_848 = _RAND_848[255:0];
  _RAND_849 = {8{`RANDOM}};
  mem_849 = _RAND_849[255:0];
  _RAND_850 = {8{`RANDOM}};
  mem_850 = _RAND_850[255:0];
  _RAND_851 = {8{`RANDOM}};
  mem_851 = _RAND_851[255:0];
  _RAND_852 = {8{`RANDOM}};
  mem_852 = _RAND_852[255:0];
  _RAND_853 = {8{`RANDOM}};
  mem_853 = _RAND_853[255:0];
  _RAND_854 = {8{`RANDOM}};
  mem_854 = _RAND_854[255:0];
  _RAND_855 = {8{`RANDOM}};
  mem_855 = _RAND_855[255:0];
  _RAND_856 = {8{`RANDOM}};
  mem_856 = _RAND_856[255:0];
  _RAND_857 = {8{`RANDOM}};
  mem_857 = _RAND_857[255:0];
  _RAND_858 = {8{`RANDOM}};
  mem_858 = _RAND_858[255:0];
  _RAND_859 = {8{`RANDOM}};
  mem_859 = _RAND_859[255:0];
  _RAND_860 = {8{`RANDOM}};
  mem_860 = _RAND_860[255:0];
  _RAND_861 = {8{`RANDOM}};
  mem_861 = _RAND_861[255:0];
  _RAND_862 = {8{`RANDOM}};
  mem_862 = _RAND_862[255:0];
  _RAND_863 = {8{`RANDOM}};
  mem_863 = _RAND_863[255:0];
  _RAND_864 = {8{`RANDOM}};
  mem_864 = _RAND_864[255:0];
  _RAND_865 = {8{`RANDOM}};
  mem_865 = _RAND_865[255:0];
  _RAND_866 = {8{`RANDOM}};
  mem_866 = _RAND_866[255:0];
  _RAND_867 = {8{`RANDOM}};
  mem_867 = _RAND_867[255:0];
  _RAND_868 = {8{`RANDOM}};
  mem_868 = _RAND_868[255:0];
  _RAND_869 = {8{`RANDOM}};
  mem_869 = _RAND_869[255:0];
  _RAND_870 = {8{`RANDOM}};
  mem_870 = _RAND_870[255:0];
  _RAND_871 = {8{`RANDOM}};
  mem_871 = _RAND_871[255:0];
  _RAND_872 = {8{`RANDOM}};
  mem_872 = _RAND_872[255:0];
  _RAND_873 = {8{`RANDOM}};
  mem_873 = _RAND_873[255:0];
  _RAND_874 = {8{`RANDOM}};
  mem_874 = _RAND_874[255:0];
  _RAND_875 = {8{`RANDOM}};
  mem_875 = _RAND_875[255:0];
  _RAND_876 = {8{`RANDOM}};
  mem_876 = _RAND_876[255:0];
  _RAND_877 = {8{`RANDOM}};
  mem_877 = _RAND_877[255:0];
  _RAND_878 = {8{`RANDOM}};
  mem_878 = _RAND_878[255:0];
  _RAND_879 = {8{`RANDOM}};
  mem_879 = _RAND_879[255:0];
  _RAND_880 = {8{`RANDOM}};
  mem_880 = _RAND_880[255:0];
  _RAND_881 = {8{`RANDOM}};
  mem_881 = _RAND_881[255:0];
  _RAND_882 = {8{`RANDOM}};
  mem_882 = _RAND_882[255:0];
  _RAND_883 = {8{`RANDOM}};
  mem_883 = _RAND_883[255:0];
  _RAND_884 = {8{`RANDOM}};
  mem_884 = _RAND_884[255:0];
  _RAND_885 = {8{`RANDOM}};
  mem_885 = _RAND_885[255:0];
  _RAND_886 = {8{`RANDOM}};
  mem_886 = _RAND_886[255:0];
  _RAND_887 = {8{`RANDOM}};
  mem_887 = _RAND_887[255:0];
  _RAND_888 = {8{`RANDOM}};
  mem_888 = _RAND_888[255:0];
  _RAND_889 = {8{`RANDOM}};
  mem_889 = _RAND_889[255:0];
  _RAND_890 = {8{`RANDOM}};
  mem_890 = _RAND_890[255:0];
  _RAND_891 = {8{`RANDOM}};
  mem_891 = _RAND_891[255:0];
  _RAND_892 = {8{`RANDOM}};
  mem_892 = _RAND_892[255:0];
  _RAND_893 = {8{`RANDOM}};
  mem_893 = _RAND_893[255:0];
  _RAND_894 = {8{`RANDOM}};
  mem_894 = _RAND_894[255:0];
  _RAND_895 = {8{`RANDOM}};
  mem_895 = _RAND_895[255:0];
  _RAND_896 = {8{`RANDOM}};
  mem_896 = _RAND_896[255:0];
  _RAND_897 = {8{`RANDOM}};
  mem_897 = _RAND_897[255:0];
  _RAND_898 = {8{`RANDOM}};
  mem_898 = _RAND_898[255:0];
  _RAND_899 = {8{`RANDOM}};
  mem_899 = _RAND_899[255:0];
  _RAND_900 = {8{`RANDOM}};
  mem_900 = _RAND_900[255:0];
  _RAND_901 = {8{`RANDOM}};
  mem_901 = _RAND_901[255:0];
  _RAND_902 = {8{`RANDOM}};
  mem_902 = _RAND_902[255:0];
  _RAND_903 = {8{`RANDOM}};
  mem_903 = _RAND_903[255:0];
  _RAND_904 = {8{`RANDOM}};
  mem_904 = _RAND_904[255:0];
  _RAND_905 = {8{`RANDOM}};
  mem_905 = _RAND_905[255:0];
  _RAND_906 = {8{`RANDOM}};
  mem_906 = _RAND_906[255:0];
  _RAND_907 = {8{`RANDOM}};
  mem_907 = _RAND_907[255:0];
  _RAND_908 = {8{`RANDOM}};
  mem_908 = _RAND_908[255:0];
  _RAND_909 = {8{`RANDOM}};
  mem_909 = _RAND_909[255:0];
  _RAND_910 = {8{`RANDOM}};
  mem_910 = _RAND_910[255:0];
  _RAND_911 = {8{`RANDOM}};
  mem_911 = _RAND_911[255:0];
  _RAND_912 = {8{`RANDOM}};
  mem_912 = _RAND_912[255:0];
  _RAND_913 = {8{`RANDOM}};
  mem_913 = _RAND_913[255:0];
  _RAND_914 = {8{`RANDOM}};
  mem_914 = _RAND_914[255:0];
  _RAND_915 = {8{`RANDOM}};
  mem_915 = _RAND_915[255:0];
  _RAND_916 = {8{`RANDOM}};
  mem_916 = _RAND_916[255:0];
  _RAND_917 = {8{`RANDOM}};
  mem_917 = _RAND_917[255:0];
  _RAND_918 = {8{`RANDOM}};
  mem_918 = _RAND_918[255:0];
  _RAND_919 = {8{`RANDOM}};
  mem_919 = _RAND_919[255:0];
  _RAND_920 = {8{`RANDOM}};
  mem_920 = _RAND_920[255:0];
  _RAND_921 = {8{`RANDOM}};
  mem_921 = _RAND_921[255:0];
  _RAND_922 = {8{`RANDOM}};
  mem_922 = _RAND_922[255:0];
  _RAND_923 = {8{`RANDOM}};
  mem_923 = _RAND_923[255:0];
  _RAND_924 = {8{`RANDOM}};
  mem_924 = _RAND_924[255:0];
  _RAND_925 = {8{`RANDOM}};
  mem_925 = _RAND_925[255:0];
  _RAND_926 = {8{`RANDOM}};
  mem_926 = _RAND_926[255:0];
  _RAND_927 = {8{`RANDOM}};
  mem_927 = _RAND_927[255:0];
  _RAND_928 = {8{`RANDOM}};
  mem_928 = _RAND_928[255:0];
  _RAND_929 = {8{`RANDOM}};
  mem_929 = _RAND_929[255:0];
  _RAND_930 = {8{`RANDOM}};
  mem_930 = _RAND_930[255:0];
  _RAND_931 = {8{`RANDOM}};
  mem_931 = _RAND_931[255:0];
  _RAND_932 = {8{`RANDOM}};
  mem_932 = _RAND_932[255:0];
  _RAND_933 = {8{`RANDOM}};
  mem_933 = _RAND_933[255:0];
  _RAND_934 = {8{`RANDOM}};
  mem_934 = _RAND_934[255:0];
  _RAND_935 = {8{`RANDOM}};
  mem_935 = _RAND_935[255:0];
  _RAND_936 = {8{`RANDOM}};
  mem_936 = _RAND_936[255:0];
  _RAND_937 = {8{`RANDOM}};
  mem_937 = _RAND_937[255:0];
  _RAND_938 = {8{`RANDOM}};
  mem_938 = _RAND_938[255:0];
  _RAND_939 = {8{`RANDOM}};
  mem_939 = _RAND_939[255:0];
  _RAND_940 = {8{`RANDOM}};
  mem_940 = _RAND_940[255:0];
  _RAND_941 = {8{`RANDOM}};
  mem_941 = _RAND_941[255:0];
  _RAND_942 = {8{`RANDOM}};
  mem_942 = _RAND_942[255:0];
  _RAND_943 = {8{`RANDOM}};
  mem_943 = _RAND_943[255:0];
  _RAND_944 = {8{`RANDOM}};
  mem_944 = _RAND_944[255:0];
  _RAND_945 = {8{`RANDOM}};
  mem_945 = _RAND_945[255:0];
  _RAND_946 = {8{`RANDOM}};
  mem_946 = _RAND_946[255:0];
  _RAND_947 = {8{`RANDOM}};
  mem_947 = _RAND_947[255:0];
  _RAND_948 = {8{`RANDOM}};
  mem_948 = _RAND_948[255:0];
  _RAND_949 = {8{`RANDOM}};
  mem_949 = _RAND_949[255:0];
  _RAND_950 = {8{`RANDOM}};
  mem_950 = _RAND_950[255:0];
  _RAND_951 = {8{`RANDOM}};
  mem_951 = _RAND_951[255:0];
  _RAND_952 = {8{`RANDOM}};
  mem_952 = _RAND_952[255:0];
  _RAND_953 = {8{`RANDOM}};
  mem_953 = _RAND_953[255:0];
  _RAND_954 = {8{`RANDOM}};
  mem_954 = _RAND_954[255:0];
  _RAND_955 = {8{`RANDOM}};
  mem_955 = _RAND_955[255:0];
  _RAND_956 = {8{`RANDOM}};
  mem_956 = _RAND_956[255:0];
  _RAND_957 = {8{`RANDOM}};
  mem_957 = _RAND_957[255:0];
  _RAND_958 = {8{`RANDOM}};
  mem_958 = _RAND_958[255:0];
  _RAND_959 = {8{`RANDOM}};
  mem_959 = _RAND_959[255:0];
  _RAND_960 = {8{`RANDOM}};
  mem_960 = _RAND_960[255:0];
  _RAND_961 = {8{`RANDOM}};
  mem_961 = _RAND_961[255:0];
  _RAND_962 = {8{`RANDOM}};
  mem_962 = _RAND_962[255:0];
  _RAND_963 = {8{`RANDOM}};
  mem_963 = _RAND_963[255:0];
  _RAND_964 = {8{`RANDOM}};
  mem_964 = _RAND_964[255:0];
  _RAND_965 = {8{`RANDOM}};
  mem_965 = _RAND_965[255:0];
  _RAND_966 = {8{`RANDOM}};
  mem_966 = _RAND_966[255:0];
  _RAND_967 = {8{`RANDOM}};
  mem_967 = _RAND_967[255:0];
  _RAND_968 = {8{`RANDOM}};
  mem_968 = _RAND_968[255:0];
  _RAND_969 = {8{`RANDOM}};
  mem_969 = _RAND_969[255:0];
  _RAND_970 = {8{`RANDOM}};
  mem_970 = _RAND_970[255:0];
  _RAND_971 = {8{`RANDOM}};
  mem_971 = _RAND_971[255:0];
  _RAND_972 = {8{`RANDOM}};
  mem_972 = _RAND_972[255:0];
  _RAND_973 = {8{`RANDOM}};
  mem_973 = _RAND_973[255:0];
  _RAND_974 = {8{`RANDOM}};
  mem_974 = _RAND_974[255:0];
  _RAND_975 = {8{`RANDOM}};
  mem_975 = _RAND_975[255:0];
  _RAND_976 = {8{`RANDOM}};
  mem_976 = _RAND_976[255:0];
  _RAND_977 = {8{`RANDOM}};
  mem_977 = _RAND_977[255:0];
  _RAND_978 = {8{`RANDOM}};
  mem_978 = _RAND_978[255:0];
  _RAND_979 = {8{`RANDOM}};
  mem_979 = _RAND_979[255:0];
  _RAND_980 = {8{`RANDOM}};
  mem_980 = _RAND_980[255:0];
  _RAND_981 = {8{`RANDOM}};
  mem_981 = _RAND_981[255:0];
  _RAND_982 = {8{`RANDOM}};
  mem_982 = _RAND_982[255:0];
  _RAND_983 = {8{`RANDOM}};
  mem_983 = _RAND_983[255:0];
  _RAND_984 = {8{`RANDOM}};
  mem_984 = _RAND_984[255:0];
  _RAND_985 = {8{`RANDOM}};
  mem_985 = _RAND_985[255:0];
  _RAND_986 = {8{`RANDOM}};
  mem_986 = _RAND_986[255:0];
  _RAND_987 = {8{`RANDOM}};
  mem_987 = _RAND_987[255:0];
  _RAND_988 = {8{`RANDOM}};
  mem_988 = _RAND_988[255:0];
  _RAND_989 = {8{`RANDOM}};
  mem_989 = _RAND_989[255:0];
  _RAND_990 = {8{`RANDOM}};
  mem_990 = _RAND_990[255:0];
  _RAND_991 = {8{`RANDOM}};
  mem_991 = _RAND_991[255:0];
  _RAND_992 = {8{`RANDOM}};
  mem_992 = _RAND_992[255:0];
  _RAND_993 = {8{`RANDOM}};
  mem_993 = _RAND_993[255:0];
  _RAND_994 = {8{`RANDOM}};
  mem_994 = _RAND_994[255:0];
  _RAND_995 = {8{`RANDOM}};
  mem_995 = _RAND_995[255:0];
  _RAND_996 = {8{`RANDOM}};
  mem_996 = _RAND_996[255:0];
  _RAND_997 = {8{`RANDOM}};
  mem_997 = _RAND_997[255:0];
  _RAND_998 = {8{`RANDOM}};
  mem_998 = _RAND_998[255:0];
  _RAND_999 = {8{`RANDOM}};
  mem_999 = _RAND_999[255:0];
  _RAND_1000 = {8{`RANDOM}};
  mem_1000 = _RAND_1000[255:0];
  _RAND_1001 = {8{`RANDOM}};
  mem_1001 = _RAND_1001[255:0];
  _RAND_1002 = {8{`RANDOM}};
  mem_1002 = _RAND_1002[255:0];
  _RAND_1003 = {8{`RANDOM}};
  mem_1003 = _RAND_1003[255:0];
  _RAND_1004 = {8{`RANDOM}};
  mem_1004 = _RAND_1004[255:0];
  _RAND_1005 = {8{`RANDOM}};
  mem_1005 = _RAND_1005[255:0];
  _RAND_1006 = {8{`RANDOM}};
  mem_1006 = _RAND_1006[255:0];
  _RAND_1007 = {8{`RANDOM}};
  mem_1007 = _RAND_1007[255:0];
  _RAND_1008 = {8{`RANDOM}};
  mem_1008 = _RAND_1008[255:0];
  _RAND_1009 = {8{`RANDOM}};
  mem_1009 = _RAND_1009[255:0];
  _RAND_1010 = {8{`RANDOM}};
  mem_1010 = _RAND_1010[255:0];
  _RAND_1011 = {8{`RANDOM}};
  mem_1011 = _RAND_1011[255:0];
  _RAND_1012 = {8{`RANDOM}};
  mem_1012 = _RAND_1012[255:0];
  _RAND_1013 = {8{`RANDOM}};
  mem_1013 = _RAND_1013[255:0];
  _RAND_1014 = {8{`RANDOM}};
  mem_1014 = _RAND_1014[255:0];
  _RAND_1015 = {8{`RANDOM}};
  mem_1015 = _RAND_1015[255:0];
  _RAND_1016 = {8{`RANDOM}};
  mem_1016 = _RAND_1016[255:0];
  _RAND_1017 = {8{`RANDOM}};
  mem_1017 = _RAND_1017[255:0];
  _RAND_1018 = {8{`RANDOM}};
  mem_1018 = _RAND_1018[255:0];
  _RAND_1019 = {8{`RANDOM}};
  mem_1019 = _RAND_1019[255:0];
  _RAND_1020 = {8{`RANDOM}};
  mem_1020 = _RAND_1020[255:0];
  _RAND_1021 = {8{`RANDOM}};
  mem_1021 = _RAND_1021[255:0];
  _RAND_1022 = {8{`RANDOM}};
  mem_1022 = _RAND_1022[255:0];
  _RAND_1023 = {8{`RANDOM}};
  mem_1023 = _RAND_1023[255:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
