module CAMLine(
  input          clock,
  input          io_we,
  input          io_wi,
  input  [127:0] io_key,
  input  [127:0] io_din,
  output         io_hit
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  write = io_we & io_wi; // @[cam.scala 58:18]
  reg [127:0] camCells; // @[cam.scala 59:21]
  assign io_hit = camCells == io_key; // @[cam.scala 65:23]
  always @(posedge clock) begin
    if (write) begin // @[cam.scala 61:14]
      camCells <= io_din; // @[cam.scala 62:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  camCells = _RAND_0[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CAM_m_n(
  input          clock,
  input          reset,
  input          io_we,
  input  [127:0] io_key,
  input  [127:0] io_din,
  input  [127:0] io_waddr,
  output         io_hit
);
  wire  CAMLine_clock; // @[cam.scala 81:36]
  wire  CAMLine_io_we; // @[cam.scala 81:36]
  wire  CAMLine_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_io_din; // @[cam.scala 81:36]
  wire  CAMLine_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_1_clock; // @[cam.scala 81:36]
  wire  CAMLine_1_io_we; // @[cam.scala 81:36]
  wire  CAMLine_1_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_1_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_1_io_din; // @[cam.scala 81:36]
  wire  CAMLine_1_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_2_clock; // @[cam.scala 81:36]
  wire  CAMLine_2_io_we; // @[cam.scala 81:36]
  wire  CAMLine_2_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_2_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_2_io_din; // @[cam.scala 81:36]
  wire  CAMLine_2_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_3_clock; // @[cam.scala 81:36]
  wire  CAMLine_3_io_we; // @[cam.scala 81:36]
  wire  CAMLine_3_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_3_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_3_io_din; // @[cam.scala 81:36]
  wire  CAMLine_3_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_4_clock; // @[cam.scala 81:36]
  wire  CAMLine_4_io_we; // @[cam.scala 81:36]
  wire  CAMLine_4_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_4_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_4_io_din; // @[cam.scala 81:36]
  wire  CAMLine_4_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_5_clock; // @[cam.scala 81:36]
  wire  CAMLine_5_io_we; // @[cam.scala 81:36]
  wire  CAMLine_5_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_5_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_5_io_din; // @[cam.scala 81:36]
  wire  CAMLine_5_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_6_clock; // @[cam.scala 81:36]
  wire  CAMLine_6_io_we; // @[cam.scala 81:36]
  wire  CAMLine_6_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_6_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_6_io_din; // @[cam.scala 81:36]
  wire  CAMLine_6_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_7_clock; // @[cam.scala 81:36]
  wire  CAMLine_7_io_we; // @[cam.scala 81:36]
  wire  CAMLine_7_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_7_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_7_io_din; // @[cam.scala 81:36]
  wire  CAMLine_7_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_8_clock; // @[cam.scala 81:36]
  wire  CAMLine_8_io_we; // @[cam.scala 81:36]
  wire  CAMLine_8_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_8_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_8_io_din; // @[cam.scala 81:36]
  wire  CAMLine_8_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_9_clock; // @[cam.scala 81:36]
  wire  CAMLine_9_io_we; // @[cam.scala 81:36]
  wire  CAMLine_9_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_9_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_9_io_din; // @[cam.scala 81:36]
  wire  CAMLine_9_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_10_clock; // @[cam.scala 81:36]
  wire  CAMLine_10_io_we; // @[cam.scala 81:36]
  wire  CAMLine_10_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_10_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_10_io_din; // @[cam.scala 81:36]
  wire  CAMLine_10_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_11_clock; // @[cam.scala 81:36]
  wire  CAMLine_11_io_we; // @[cam.scala 81:36]
  wire  CAMLine_11_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_11_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_11_io_din; // @[cam.scala 81:36]
  wire  CAMLine_11_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_12_clock; // @[cam.scala 81:36]
  wire  CAMLine_12_io_we; // @[cam.scala 81:36]
  wire  CAMLine_12_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_12_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_12_io_din; // @[cam.scala 81:36]
  wire  CAMLine_12_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_13_clock; // @[cam.scala 81:36]
  wire  CAMLine_13_io_we; // @[cam.scala 81:36]
  wire  CAMLine_13_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_13_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_13_io_din; // @[cam.scala 81:36]
  wire  CAMLine_13_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_14_clock; // @[cam.scala 81:36]
  wire  CAMLine_14_io_we; // @[cam.scala 81:36]
  wire  CAMLine_14_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_14_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_14_io_din; // @[cam.scala 81:36]
  wire  CAMLine_14_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_15_clock; // @[cam.scala 81:36]
  wire  CAMLine_15_io_we; // @[cam.scala 81:36]
  wire  CAMLine_15_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_15_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_15_io_din; // @[cam.scala 81:36]
  wire  CAMLine_15_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_16_clock; // @[cam.scala 81:36]
  wire  CAMLine_16_io_we; // @[cam.scala 81:36]
  wire  CAMLine_16_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_16_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_16_io_din; // @[cam.scala 81:36]
  wire  CAMLine_16_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_17_clock; // @[cam.scala 81:36]
  wire  CAMLine_17_io_we; // @[cam.scala 81:36]
  wire  CAMLine_17_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_17_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_17_io_din; // @[cam.scala 81:36]
  wire  CAMLine_17_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_18_clock; // @[cam.scala 81:36]
  wire  CAMLine_18_io_we; // @[cam.scala 81:36]
  wire  CAMLine_18_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_18_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_18_io_din; // @[cam.scala 81:36]
  wire  CAMLine_18_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_19_clock; // @[cam.scala 81:36]
  wire  CAMLine_19_io_we; // @[cam.scala 81:36]
  wire  CAMLine_19_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_19_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_19_io_din; // @[cam.scala 81:36]
  wire  CAMLine_19_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_20_clock; // @[cam.scala 81:36]
  wire  CAMLine_20_io_we; // @[cam.scala 81:36]
  wire  CAMLine_20_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_20_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_20_io_din; // @[cam.scala 81:36]
  wire  CAMLine_20_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_21_clock; // @[cam.scala 81:36]
  wire  CAMLine_21_io_we; // @[cam.scala 81:36]
  wire  CAMLine_21_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_21_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_21_io_din; // @[cam.scala 81:36]
  wire  CAMLine_21_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_22_clock; // @[cam.scala 81:36]
  wire  CAMLine_22_io_we; // @[cam.scala 81:36]
  wire  CAMLine_22_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_22_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_22_io_din; // @[cam.scala 81:36]
  wire  CAMLine_22_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_23_clock; // @[cam.scala 81:36]
  wire  CAMLine_23_io_we; // @[cam.scala 81:36]
  wire  CAMLine_23_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_23_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_23_io_din; // @[cam.scala 81:36]
  wire  CAMLine_23_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_24_clock; // @[cam.scala 81:36]
  wire  CAMLine_24_io_we; // @[cam.scala 81:36]
  wire  CAMLine_24_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_24_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_24_io_din; // @[cam.scala 81:36]
  wire  CAMLine_24_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_25_clock; // @[cam.scala 81:36]
  wire  CAMLine_25_io_we; // @[cam.scala 81:36]
  wire  CAMLine_25_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_25_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_25_io_din; // @[cam.scala 81:36]
  wire  CAMLine_25_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_26_clock; // @[cam.scala 81:36]
  wire  CAMLine_26_io_we; // @[cam.scala 81:36]
  wire  CAMLine_26_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_26_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_26_io_din; // @[cam.scala 81:36]
  wire  CAMLine_26_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_27_clock; // @[cam.scala 81:36]
  wire  CAMLine_27_io_we; // @[cam.scala 81:36]
  wire  CAMLine_27_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_27_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_27_io_din; // @[cam.scala 81:36]
  wire  CAMLine_27_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_28_clock; // @[cam.scala 81:36]
  wire  CAMLine_28_io_we; // @[cam.scala 81:36]
  wire  CAMLine_28_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_28_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_28_io_din; // @[cam.scala 81:36]
  wire  CAMLine_28_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_29_clock; // @[cam.scala 81:36]
  wire  CAMLine_29_io_we; // @[cam.scala 81:36]
  wire  CAMLine_29_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_29_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_29_io_din; // @[cam.scala 81:36]
  wire  CAMLine_29_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_30_clock; // @[cam.scala 81:36]
  wire  CAMLine_30_io_we; // @[cam.scala 81:36]
  wire  CAMLine_30_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_30_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_30_io_din; // @[cam.scala 81:36]
  wire  CAMLine_30_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_31_clock; // @[cam.scala 81:36]
  wire  CAMLine_31_io_we; // @[cam.scala 81:36]
  wire  CAMLine_31_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_31_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_31_io_din; // @[cam.scala 81:36]
  wire  CAMLine_31_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_32_clock; // @[cam.scala 81:36]
  wire  CAMLine_32_io_we; // @[cam.scala 81:36]
  wire  CAMLine_32_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_32_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_32_io_din; // @[cam.scala 81:36]
  wire  CAMLine_32_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_33_clock; // @[cam.scala 81:36]
  wire  CAMLine_33_io_we; // @[cam.scala 81:36]
  wire  CAMLine_33_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_33_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_33_io_din; // @[cam.scala 81:36]
  wire  CAMLine_33_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_34_clock; // @[cam.scala 81:36]
  wire  CAMLine_34_io_we; // @[cam.scala 81:36]
  wire  CAMLine_34_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_34_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_34_io_din; // @[cam.scala 81:36]
  wire  CAMLine_34_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_35_clock; // @[cam.scala 81:36]
  wire  CAMLine_35_io_we; // @[cam.scala 81:36]
  wire  CAMLine_35_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_35_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_35_io_din; // @[cam.scala 81:36]
  wire  CAMLine_35_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_36_clock; // @[cam.scala 81:36]
  wire  CAMLine_36_io_we; // @[cam.scala 81:36]
  wire  CAMLine_36_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_36_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_36_io_din; // @[cam.scala 81:36]
  wire  CAMLine_36_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_37_clock; // @[cam.scala 81:36]
  wire  CAMLine_37_io_we; // @[cam.scala 81:36]
  wire  CAMLine_37_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_37_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_37_io_din; // @[cam.scala 81:36]
  wire  CAMLine_37_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_38_clock; // @[cam.scala 81:36]
  wire  CAMLine_38_io_we; // @[cam.scala 81:36]
  wire  CAMLine_38_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_38_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_38_io_din; // @[cam.scala 81:36]
  wire  CAMLine_38_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_39_clock; // @[cam.scala 81:36]
  wire  CAMLine_39_io_we; // @[cam.scala 81:36]
  wire  CAMLine_39_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_39_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_39_io_din; // @[cam.scala 81:36]
  wire  CAMLine_39_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_40_clock; // @[cam.scala 81:36]
  wire  CAMLine_40_io_we; // @[cam.scala 81:36]
  wire  CAMLine_40_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_40_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_40_io_din; // @[cam.scala 81:36]
  wire  CAMLine_40_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_41_clock; // @[cam.scala 81:36]
  wire  CAMLine_41_io_we; // @[cam.scala 81:36]
  wire  CAMLine_41_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_41_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_41_io_din; // @[cam.scala 81:36]
  wire  CAMLine_41_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_42_clock; // @[cam.scala 81:36]
  wire  CAMLine_42_io_we; // @[cam.scala 81:36]
  wire  CAMLine_42_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_42_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_42_io_din; // @[cam.scala 81:36]
  wire  CAMLine_42_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_43_clock; // @[cam.scala 81:36]
  wire  CAMLine_43_io_we; // @[cam.scala 81:36]
  wire  CAMLine_43_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_43_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_43_io_din; // @[cam.scala 81:36]
  wire  CAMLine_43_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_44_clock; // @[cam.scala 81:36]
  wire  CAMLine_44_io_we; // @[cam.scala 81:36]
  wire  CAMLine_44_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_44_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_44_io_din; // @[cam.scala 81:36]
  wire  CAMLine_44_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_45_clock; // @[cam.scala 81:36]
  wire  CAMLine_45_io_we; // @[cam.scala 81:36]
  wire  CAMLine_45_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_45_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_45_io_din; // @[cam.scala 81:36]
  wire  CAMLine_45_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_46_clock; // @[cam.scala 81:36]
  wire  CAMLine_46_io_we; // @[cam.scala 81:36]
  wire  CAMLine_46_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_46_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_46_io_din; // @[cam.scala 81:36]
  wire  CAMLine_46_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_47_clock; // @[cam.scala 81:36]
  wire  CAMLine_47_io_we; // @[cam.scala 81:36]
  wire  CAMLine_47_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_47_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_47_io_din; // @[cam.scala 81:36]
  wire  CAMLine_47_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_48_clock; // @[cam.scala 81:36]
  wire  CAMLine_48_io_we; // @[cam.scala 81:36]
  wire  CAMLine_48_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_48_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_48_io_din; // @[cam.scala 81:36]
  wire  CAMLine_48_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_49_clock; // @[cam.scala 81:36]
  wire  CAMLine_49_io_we; // @[cam.scala 81:36]
  wire  CAMLine_49_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_49_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_49_io_din; // @[cam.scala 81:36]
  wire  CAMLine_49_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_50_clock; // @[cam.scala 81:36]
  wire  CAMLine_50_io_we; // @[cam.scala 81:36]
  wire  CAMLine_50_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_50_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_50_io_din; // @[cam.scala 81:36]
  wire  CAMLine_50_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_51_clock; // @[cam.scala 81:36]
  wire  CAMLine_51_io_we; // @[cam.scala 81:36]
  wire  CAMLine_51_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_51_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_51_io_din; // @[cam.scala 81:36]
  wire  CAMLine_51_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_52_clock; // @[cam.scala 81:36]
  wire  CAMLine_52_io_we; // @[cam.scala 81:36]
  wire  CAMLine_52_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_52_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_52_io_din; // @[cam.scala 81:36]
  wire  CAMLine_52_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_53_clock; // @[cam.scala 81:36]
  wire  CAMLine_53_io_we; // @[cam.scala 81:36]
  wire  CAMLine_53_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_53_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_53_io_din; // @[cam.scala 81:36]
  wire  CAMLine_53_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_54_clock; // @[cam.scala 81:36]
  wire  CAMLine_54_io_we; // @[cam.scala 81:36]
  wire  CAMLine_54_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_54_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_54_io_din; // @[cam.scala 81:36]
  wire  CAMLine_54_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_55_clock; // @[cam.scala 81:36]
  wire  CAMLine_55_io_we; // @[cam.scala 81:36]
  wire  CAMLine_55_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_55_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_55_io_din; // @[cam.scala 81:36]
  wire  CAMLine_55_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_56_clock; // @[cam.scala 81:36]
  wire  CAMLine_56_io_we; // @[cam.scala 81:36]
  wire  CAMLine_56_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_56_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_56_io_din; // @[cam.scala 81:36]
  wire  CAMLine_56_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_57_clock; // @[cam.scala 81:36]
  wire  CAMLine_57_io_we; // @[cam.scala 81:36]
  wire  CAMLine_57_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_57_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_57_io_din; // @[cam.scala 81:36]
  wire  CAMLine_57_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_58_clock; // @[cam.scala 81:36]
  wire  CAMLine_58_io_we; // @[cam.scala 81:36]
  wire  CAMLine_58_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_58_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_58_io_din; // @[cam.scala 81:36]
  wire  CAMLine_58_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_59_clock; // @[cam.scala 81:36]
  wire  CAMLine_59_io_we; // @[cam.scala 81:36]
  wire  CAMLine_59_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_59_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_59_io_din; // @[cam.scala 81:36]
  wire  CAMLine_59_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_60_clock; // @[cam.scala 81:36]
  wire  CAMLine_60_io_we; // @[cam.scala 81:36]
  wire  CAMLine_60_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_60_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_60_io_din; // @[cam.scala 81:36]
  wire  CAMLine_60_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_61_clock; // @[cam.scala 81:36]
  wire  CAMLine_61_io_we; // @[cam.scala 81:36]
  wire  CAMLine_61_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_61_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_61_io_din; // @[cam.scala 81:36]
  wire  CAMLine_61_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_62_clock; // @[cam.scala 81:36]
  wire  CAMLine_62_io_we; // @[cam.scala 81:36]
  wire  CAMLine_62_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_62_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_62_io_din; // @[cam.scala 81:36]
  wire  CAMLine_62_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_63_clock; // @[cam.scala 81:36]
  wire  CAMLine_63_io_we; // @[cam.scala 81:36]
  wire  CAMLine_63_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_63_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_63_io_din; // @[cam.scala 81:36]
  wire  CAMLine_63_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_64_clock; // @[cam.scala 81:36]
  wire  CAMLine_64_io_we; // @[cam.scala 81:36]
  wire  CAMLine_64_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_64_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_64_io_din; // @[cam.scala 81:36]
  wire  CAMLine_64_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_65_clock; // @[cam.scala 81:36]
  wire  CAMLine_65_io_we; // @[cam.scala 81:36]
  wire  CAMLine_65_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_65_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_65_io_din; // @[cam.scala 81:36]
  wire  CAMLine_65_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_66_clock; // @[cam.scala 81:36]
  wire  CAMLine_66_io_we; // @[cam.scala 81:36]
  wire  CAMLine_66_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_66_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_66_io_din; // @[cam.scala 81:36]
  wire  CAMLine_66_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_67_clock; // @[cam.scala 81:36]
  wire  CAMLine_67_io_we; // @[cam.scala 81:36]
  wire  CAMLine_67_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_67_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_67_io_din; // @[cam.scala 81:36]
  wire  CAMLine_67_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_68_clock; // @[cam.scala 81:36]
  wire  CAMLine_68_io_we; // @[cam.scala 81:36]
  wire  CAMLine_68_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_68_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_68_io_din; // @[cam.scala 81:36]
  wire  CAMLine_68_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_69_clock; // @[cam.scala 81:36]
  wire  CAMLine_69_io_we; // @[cam.scala 81:36]
  wire  CAMLine_69_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_69_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_69_io_din; // @[cam.scala 81:36]
  wire  CAMLine_69_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_70_clock; // @[cam.scala 81:36]
  wire  CAMLine_70_io_we; // @[cam.scala 81:36]
  wire  CAMLine_70_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_70_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_70_io_din; // @[cam.scala 81:36]
  wire  CAMLine_70_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_71_clock; // @[cam.scala 81:36]
  wire  CAMLine_71_io_we; // @[cam.scala 81:36]
  wire  CAMLine_71_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_71_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_71_io_din; // @[cam.scala 81:36]
  wire  CAMLine_71_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_72_clock; // @[cam.scala 81:36]
  wire  CAMLine_72_io_we; // @[cam.scala 81:36]
  wire  CAMLine_72_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_72_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_72_io_din; // @[cam.scala 81:36]
  wire  CAMLine_72_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_73_clock; // @[cam.scala 81:36]
  wire  CAMLine_73_io_we; // @[cam.scala 81:36]
  wire  CAMLine_73_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_73_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_73_io_din; // @[cam.scala 81:36]
  wire  CAMLine_73_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_74_clock; // @[cam.scala 81:36]
  wire  CAMLine_74_io_we; // @[cam.scala 81:36]
  wire  CAMLine_74_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_74_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_74_io_din; // @[cam.scala 81:36]
  wire  CAMLine_74_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_75_clock; // @[cam.scala 81:36]
  wire  CAMLine_75_io_we; // @[cam.scala 81:36]
  wire  CAMLine_75_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_75_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_75_io_din; // @[cam.scala 81:36]
  wire  CAMLine_75_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_76_clock; // @[cam.scala 81:36]
  wire  CAMLine_76_io_we; // @[cam.scala 81:36]
  wire  CAMLine_76_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_76_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_76_io_din; // @[cam.scala 81:36]
  wire  CAMLine_76_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_77_clock; // @[cam.scala 81:36]
  wire  CAMLine_77_io_we; // @[cam.scala 81:36]
  wire  CAMLine_77_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_77_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_77_io_din; // @[cam.scala 81:36]
  wire  CAMLine_77_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_78_clock; // @[cam.scala 81:36]
  wire  CAMLine_78_io_we; // @[cam.scala 81:36]
  wire  CAMLine_78_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_78_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_78_io_din; // @[cam.scala 81:36]
  wire  CAMLine_78_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_79_clock; // @[cam.scala 81:36]
  wire  CAMLine_79_io_we; // @[cam.scala 81:36]
  wire  CAMLine_79_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_79_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_79_io_din; // @[cam.scala 81:36]
  wire  CAMLine_79_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_80_clock; // @[cam.scala 81:36]
  wire  CAMLine_80_io_we; // @[cam.scala 81:36]
  wire  CAMLine_80_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_80_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_80_io_din; // @[cam.scala 81:36]
  wire  CAMLine_80_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_81_clock; // @[cam.scala 81:36]
  wire  CAMLine_81_io_we; // @[cam.scala 81:36]
  wire  CAMLine_81_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_81_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_81_io_din; // @[cam.scala 81:36]
  wire  CAMLine_81_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_82_clock; // @[cam.scala 81:36]
  wire  CAMLine_82_io_we; // @[cam.scala 81:36]
  wire  CAMLine_82_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_82_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_82_io_din; // @[cam.scala 81:36]
  wire  CAMLine_82_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_83_clock; // @[cam.scala 81:36]
  wire  CAMLine_83_io_we; // @[cam.scala 81:36]
  wire  CAMLine_83_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_83_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_83_io_din; // @[cam.scala 81:36]
  wire  CAMLine_83_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_84_clock; // @[cam.scala 81:36]
  wire  CAMLine_84_io_we; // @[cam.scala 81:36]
  wire  CAMLine_84_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_84_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_84_io_din; // @[cam.scala 81:36]
  wire  CAMLine_84_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_85_clock; // @[cam.scala 81:36]
  wire  CAMLine_85_io_we; // @[cam.scala 81:36]
  wire  CAMLine_85_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_85_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_85_io_din; // @[cam.scala 81:36]
  wire  CAMLine_85_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_86_clock; // @[cam.scala 81:36]
  wire  CAMLine_86_io_we; // @[cam.scala 81:36]
  wire  CAMLine_86_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_86_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_86_io_din; // @[cam.scala 81:36]
  wire  CAMLine_86_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_87_clock; // @[cam.scala 81:36]
  wire  CAMLine_87_io_we; // @[cam.scala 81:36]
  wire  CAMLine_87_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_87_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_87_io_din; // @[cam.scala 81:36]
  wire  CAMLine_87_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_88_clock; // @[cam.scala 81:36]
  wire  CAMLine_88_io_we; // @[cam.scala 81:36]
  wire  CAMLine_88_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_88_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_88_io_din; // @[cam.scala 81:36]
  wire  CAMLine_88_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_89_clock; // @[cam.scala 81:36]
  wire  CAMLine_89_io_we; // @[cam.scala 81:36]
  wire  CAMLine_89_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_89_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_89_io_din; // @[cam.scala 81:36]
  wire  CAMLine_89_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_90_clock; // @[cam.scala 81:36]
  wire  CAMLine_90_io_we; // @[cam.scala 81:36]
  wire  CAMLine_90_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_90_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_90_io_din; // @[cam.scala 81:36]
  wire  CAMLine_90_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_91_clock; // @[cam.scala 81:36]
  wire  CAMLine_91_io_we; // @[cam.scala 81:36]
  wire  CAMLine_91_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_91_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_91_io_din; // @[cam.scala 81:36]
  wire  CAMLine_91_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_92_clock; // @[cam.scala 81:36]
  wire  CAMLine_92_io_we; // @[cam.scala 81:36]
  wire  CAMLine_92_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_92_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_92_io_din; // @[cam.scala 81:36]
  wire  CAMLine_92_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_93_clock; // @[cam.scala 81:36]
  wire  CAMLine_93_io_we; // @[cam.scala 81:36]
  wire  CAMLine_93_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_93_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_93_io_din; // @[cam.scala 81:36]
  wire  CAMLine_93_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_94_clock; // @[cam.scala 81:36]
  wire  CAMLine_94_io_we; // @[cam.scala 81:36]
  wire  CAMLine_94_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_94_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_94_io_din; // @[cam.scala 81:36]
  wire  CAMLine_94_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_95_clock; // @[cam.scala 81:36]
  wire  CAMLine_95_io_we; // @[cam.scala 81:36]
  wire  CAMLine_95_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_95_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_95_io_din; // @[cam.scala 81:36]
  wire  CAMLine_95_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_96_clock; // @[cam.scala 81:36]
  wire  CAMLine_96_io_we; // @[cam.scala 81:36]
  wire  CAMLine_96_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_96_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_96_io_din; // @[cam.scala 81:36]
  wire  CAMLine_96_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_97_clock; // @[cam.scala 81:36]
  wire  CAMLine_97_io_we; // @[cam.scala 81:36]
  wire  CAMLine_97_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_97_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_97_io_din; // @[cam.scala 81:36]
  wire  CAMLine_97_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_98_clock; // @[cam.scala 81:36]
  wire  CAMLine_98_io_we; // @[cam.scala 81:36]
  wire  CAMLine_98_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_98_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_98_io_din; // @[cam.scala 81:36]
  wire  CAMLine_98_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_99_clock; // @[cam.scala 81:36]
  wire  CAMLine_99_io_we; // @[cam.scala 81:36]
  wire  CAMLine_99_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_99_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_99_io_din; // @[cam.scala 81:36]
  wire  CAMLine_99_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_100_clock; // @[cam.scala 81:36]
  wire  CAMLine_100_io_we; // @[cam.scala 81:36]
  wire  CAMLine_100_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_100_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_100_io_din; // @[cam.scala 81:36]
  wire  CAMLine_100_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_101_clock; // @[cam.scala 81:36]
  wire  CAMLine_101_io_we; // @[cam.scala 81:36]
  wire  CAMLine_101_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_101_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_101_io_din; // @[cam.scala 81:36]
  wire  CAMLine_101_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_102_clock; // @[cam.scala 81:36]
  wire  CAMLine_102_io_we; // @[cam.scala 81:36]
  wire  CAMLine_102_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_102_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_102_io_din; // @[cam.scala 81:36]
  wire  CAMLine_102_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_103_clock; // @[cam.scala 81:36]
  wire  CAMLine_103_io_we; // @[cam.scala 81:36]
  wire  CAMLine_103_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_103_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_103_io_din; // @[cam.scala 81:36]
  wire  CAMLine_103_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_104_clock; // @[cam.scala 81:36]
  wire  CAMLine_104_io_we; // @[cam.scala 81:36]
  wire  CAMLine_104_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_104_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_104_io_din; // @[cam.scala 81:36]
  wire  CAMLine_104_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_105_clock; // @[cam.scala 81:36]
  wire  CAMLine_105_io_we; // @[cam.scala 81:36]
  wire  CAMLine_105_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_105_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_105_io_din; // @[cam.scala 81:36]
  wire  CAMLine_105_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_106_clock; // @[cam.scala 81:36]
  wire  CAMLine_106_io_we; // @[cam.scala 81:36]
  wire  CAMLine_106_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_106_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_106_io_din; // @[cam.scala 81:36]
  wire  CAMLine_106_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_107_clock; // @[cam.scala 81:36]
  wire  CAMLine_107_io_we; // @[cam.scala 81:36]
  wire  CAMLine_107_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_107_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_107_io_din; // @[cam.scala 81:36]
  wire  CAMLine_107_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_108_clock; // @[cam.scala 81:36]
  wire  CAMLine_108_io_we; // @[cam.scala 81:36]
  wire  CAMLine_108_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_108_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_108_io_din; // @[cam.scala 81:36]
  wire  CAMLine_108_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_109_clock; // @[cam.scala 81:36]
  wire  CAMLine_109_io_we; // @[cam.scala 81:36]
  wire  CAMLine_109_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_109_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_109_io_din; // @[cam.scala 81:36]
  wire  CAMLine_109_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_110_clock; // @[cam.scala 81:36]
  wire  CAMLine_110_io_we; // @[cam.scala 81:36]
  wire  CAMLine_110_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_110_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_110_io_din; // @[cam.scala 81:36]
  wire  CAMLine_110_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_111_clock; // @[cam.scala 81:36]
  wire  CAMLine_111_io_we; // @[cam.scala 81:36]
  wire  CAMLine_111_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_111_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_111_io_din; // @[cam.scala 81:36]
  wire  CAMLine_111_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_112_clock; // @[cam.scala 81:36]
  wire  CAMLine_112_io_we; // @[cam.scala 81:36]
  wire  CAMLine_112_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_112_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_112_io_din; // @[cam.scala 81:36]
  wire  CAMLine_112_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_113_clock; // @[cam.scala 81:36]
  wire  CAMLine_113_io_we; // @[cam.scala 81:36]
  wire  CAMLine_113_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_113_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_113_io_din; // @[cam.scala 81:36]
  wire  CAMLine_113_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_114_clock; // @[cam.scala 81:36]
  wire  CAMLine_114_io_we; // @[cam.scala 81:36]
  wire  CAMLine_114_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_114_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_114_io_din; // @[cam.scala 81:36]
  wire  CAMLine_114_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_115_clock; // @[cam.scala 81:36]
  wire  CAMLine_115_io_we; // @[cam.scala 81:36]
  wire  CAMLine_115_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_115_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_115_io_din; // @[cam.scala 81:36]
  wire  CAMLine_115_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_116_clock; // @[cam.scala 81:36]
  wire  CAMLine_116_io_we; // @[cam.scala 81:36]
  wire  CAMLine_116_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_116_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_116_io_din; // @[cam.scala 81:36]
  wire  CAMLine_116_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_117_clock; // @[cam.scala 81:36]
  wire  CAMLine_117_io_we; // @[cam.scala 81:36]
  wire  CAMLine_117_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_117_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_117_io_din; // @[cam.scala 81:36]
  wire  CAMLine_117_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_118_clock; // @[cam.scala 81:36]
  wire  CAMLine_118_io_we; // @[cam.scala 81:36]
  wire  CAMLine_118_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_118_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_118_io_din; // @[cam.scala 81:36]
  wire  CAMLine_118_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_119_clock; // @[cam.scala 81:36]
  wire  CAMLine_119_io_we; // @[cam.scala 81:36]
  wire  CAMLine_119_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_119_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_119_io_din; // @[cam.scala 81:36]
  wire  CAMLine_119_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_120_clock; // @[cam.scala 81:36]
  wire  CAMLine_120_io_we; // @[cam.scala 81:36]
  wire  CAMLine_120_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_120_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_120_io_din; // @[cam.scala 81:36]
  wire  CAMLine_120_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_121_clock; // @[cam.scala 81:36]
  wire  CAMLine_121_io_we; // @[cam.scala 81:36]
  wire  CAMLine_121_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_121_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_121_io_din; // @[cam.scala 81:36]
  wire  CAMLine_121_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_122_clock; // @[cam.scala 81:36]
  wire  CAMLine_122_io_we; // @[cam.scala 81:36]
  wire  CAMLine_122_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_122_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_122_io_din; // @[cam.scala 81:36]
  wire  CAMLine_122_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_123_clock; // @[cam.scala 81:36]
  wire  CAMLine_123_io_we; // @[cam.scala 81:36]
  wire  CAMLine_123_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_123_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_123_io_din; // @[cam.scala 81:36]
  wire  CAMLine_123_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_124_clock; // @[cam.scala 81:36]
  wire  CAMLine_124_io_we; // @[cam.scala 81:36]
  wire  CAMLine_124_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_124_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_124_io_din; // @[cam.scala 81:36]
  wire  CAMLine_124_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_125_clock; // @[cam.scala 81:36]
  wire  CAMLine_125_io_we; // @[cam.scala 81:36]
  wire  CAMLine_125_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_125_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_125_io_din; // @[cam.scala 81:36]
  wire  CAMLine_125_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_126_clock; // @[cam.scala 81:36]
  wire  CAMLine_126_io_we; // @[cam.scala 81:36]
  wire  CAMLine_126_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_126_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_126_io_din; // @[cam.scala 81:36]
  wire  CAMLine_126_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_127_clock; // @[cam.scala 81:36]
  wire  CAMLine_127_io_we; // @[cam.scala 81:36]
  wire  CAMLine_127_io_wi; // @[cam.scala 81:36]
  wire [127:0] CAMLine_127_io_key; // @[cam.scala 81:36]
  wire [127:0] CAMLine_127_io_din; // @[cam.scala 81:36]
  wire  CAMLine_127_io_hit; // @[cam.scala 81:36]
  wire  _io_hit_T_29 = CAMLine_io_hit | CAMLine_1_io_hit | CAMLine_2_io_hit | CAMLine_3_io_hit | CAMLine_4_io_hit |
    CAMLine_5_io_hit | CAMLine_6_io_hit | CAMLine_7_io_hit | CAMLine_8_io_hit | CAMLine_9_io_hit | CAMLine_10_io_hit |
    CAMLine_11_io_hit | CAMLine_12_io_hit | CAMLine_13_io_hit | CAMLine_14_io_hit | CAMLine_15_io_hit |
    CAMLine_16_io_hit | CAMLine_17_io_hit | CAMLine_18_io_hit | CAMLine_19_io_hit | CAMLine_20_io_hit |
    CAMLine_21_io_hit | CAMLine_22_io_hit | CAMLine_23_io_hit | CAMLine_24_io_hit | CAMLine_25_io_hit |
    CAMLine_26_io_hit | CAMLine_27_io_hit | CAMLine_28_io_hit | CAMLine_29_io_hit | CAMLine_30_io_hit; // @[cam.scala 93:27]
  wire  _io_hit_T_59 = _io_hit_T_29 | CAMLine_31_io_hit | CAMLine_32_io_hit | CAMLine_33_io_hit | CAMLine_34_io_hit |
    CAMLine_35_io_hit | CAMLine_36_io_hit | CAMLine_37_io_hit | CAMLine_38_io_hit | CAMLine_39_io_hit |
    CAMLine_40_io_hit | CAMLine_41_io_hit | CAMLine_42_io_hit | CAMLine_43_io_hit | CAMLine_44_io_hit |
    CAMLine_45_io_hit | CAMLine_46_io_hit | CAMLine_47_io_hit | CAMLine_48_io_hit | CAMLine_49_io_hit |
    CAMLine_50_io_hit | CAMLine_51_io_hit | CAMLine_52_io_hit | CAMLine_53_io_hit | CAMLine_54_io_hit |
    CAMLine_55_io_hit | CAMLine_56_io_hit | CAMLine_57_io_hit | CAMLine_58_io_hit | CAMLine_59_io_hit |
    CAMLine_60_io_hit; // @[cam.scala 93:27]
  wire  _io_hit_T_89 = _io_hit_T_59 | CAMLine_61_io_hit | CAMLine_62_io_hit | CAMLine_63_io_hit | CAMLine_64_io_hit |
    CAMLine_65_io_hit | CAMLine_66_io_hit | CAMLine_67_io_hit | CAMLine_68_io_hit | CAMLine_69_io_hit |
    CAMLine_70_io_hit | CAMLine_71_io_hit | CAMLine_72_io_hit | CAMLine_73_io_hit | CAMLine_74_io_hit |
    CAMLine_75_io_hit | CAMLine_76_io_hit | CAMLine_77_io_hit | CAMLine_78_io_hit | CAMLine_79_io_hit |
    CAMLine_80_io_hit | CAMLine_81_io_hit | CAMLine_82_io_hit | CAMLine_83_io_hit | CAMLine_84_io_hit |
    CAMLine_85_io_hit | CAMLine_86_io_hit | CAMLine_87_io_hit | CAMLine_88_io_hit | CAMLine_89_io_hit |
    CAMLine_90_io_hit; // @[cam.scala 93:27]
  wire  _io_hit_T_119 = _io_hit_T_89 | CAMLine_91_io_hit | CAMLine_92_io_hit | CAMLine_93_io_hit | CAMLine_94_io_hit |
    CAMLine_95_io_hit | CAMLine_96_io_hit | CAMLine_97_io_hit | CAMLine_98_io_hit | CAMLine_99_io_hit |
    CAMLine_100_io_hit | CAMLine_101_io_hit | CAMLine_102_io_hit | CAMLine_103_io_hit | CAMLine_104_io_hit |
    CAMLine_105_io_hit | CAMLine_106_io_hit | CAMLine_107_io_hit | CAMLine_108_io_hit | CAMLine_109_io_hit |
    CAMLine_110_io_hit | CAMLine_111_io_hit | CAMLine_112_io_hit | CAMLine_113_io_hit | CAMLine_114_io_hit |
    CAMLine_115_io_hit | CAMLine_116_io_hit | CAMLine_117_io_hit | CAMLine_118_io_hit | CAMLine_119_io_hit |
    CAMLine_120_io_hit; // @[cam.scala 93:27]
  CAMLine CAMLine ( // @[cam.scala 81:36]
    .clock(CAMLine_clock),
    .io_we(CAMLine_io_we),
    .io_wi(CAMLine_io_wi),
    .io_key(CAMLine_io_key),
    .io_din(CAMLine_io_din),
    .io_hit(CAMLine_io_hit)
  );
  CAMLine CAMLine_1 ( // @[cam.scala 81:36]
    .clock(CAMLine_1_clock),
    .io_we(CAMLine_1_io_we),
    .io_wi(CAMLine_1_io_wi),
    .io_key(CAMLine_1_io_key),
    .io_din(CAMLine_1_io_din),
    .io_hit(CAMLine_1_io_hit)
  );
  CAMLine CAMLine_2 ( // @[cam.scala 81:36]
    .clock(CAMLine_2_clock),
    .io_we(CAMLine_2_io_we),
    .io_wi(CAMLine_2_io_wi),
    .io_key(CAMLine_2_io_key),
    .io_din(CAMLine_2_io_din),
    .io_hit(CAMLine_2_io_hit)
  );
  CAMLine CAMLine_3 ( // @[cam.scala 81:36]
    .clock(CAMLine_3_clock),
    .io_we(CAMLine_3_io_we),
    .io_wi(CAMLine_3_io_wi),
    .io_key(CAMLine_3_io_key),
    .io_din(CAMLine_3_io_din),
    .io_hit(CAMLine_3_io_hit)
  );
  CAMLine CAMLine_4 ( // @[cam.scala 81:36]
    .clock(CAMLine_4_clock),
    .io_we(CAMLine_4_io_we),
    .io_wi(CAMLine_4_io_wi),
    .io_key(CAMLine_4_io_key),
    .io_din(CAMLine_4_io_din),
    .io_hit(CAMLine_4_io_hit)
  );
  CAMLine CAMLine_5 ( // @[cam.scala 81:36]
    .clock(CAMLine_5_clock),
    .io_we(CAMLine_5_io_we),
    .io_wi(CAMLine_5_io_wi),
    .io_key(CAMLine_5_io_key),
    .io_din(CAMLine_5_io_din),
    .io_hit(CAMLine_5_io_hit)
  );
  CAMLine CAMLine_6 ( // @[cam.scala 81:36]
    .clock(CAMLine_6_clock),
    .io_we(CAMLine_6_io_we),
    .io_wi(CAMLine_6_io_wi),
    .io_key(CAMLine_6_io_key),
    .io_din(CAMLine_6_io_din),
    .io_hit(CAMLine_6_io_hit)
  );
  CAMLine CAMLine_7 ( // @[cam.scala 81:36]
    .clock(CAMLine_7_clock),
    .io_we(CAMLine_7_io_we),
    .io_wi(CAMLine_7_io_wi),
    .io_key(CAMLine_7_io_key),
    .io_din(CAMLine_7_io_din),
    .io_hit(CAMLine_7_io_hit)
  );
  CAMLine CAMLine_8 ( // @[cam.scala 81:36]
    .clock(CAMLine_8_clock),
    .io_we(CAMLine_8_io_we),
    .io_wi(CAMLine_8_io_wi),
    .io_key(CAMLine_8_io_key),
    .io_din(CAMLine_8_io_din),
    .io_hit(CAMLine_8_io_hit)
  );
  CAMLine CAMLine_9 ( // @[cam.scala 81:36]
    .clock(CAMLine_9_clock),
    .io_we(CAMLine_9_io_we),
    .io_wi(CAMLine_9_io_wi),
    .io_key(CAMLine_9_io_key),
    .io_din(CAMLine_9_io_din),
    .io_hit(CAMLine_9_io_hit)
  );
  CAMLine CAMLine_10 ( // @[cam.scala 81:36]
    .clock(CAMLine_10_clock),
    .io_we(CAMLine_10_io_we),
    .io_wi(CAMLine_10_io_wi),
    .io_key(CAMLine_10_io_key),
    .io_din(CAMLine_10_io_din),
    .io_hit(CAMLine_10_io_hit)
  );
  CAMLine CAMLine_11 ( // @[cam.scala 81:36]
    .clock(CAMLine_11_clock),
    .io_we(CAMLine_11_io_we),
    .io_wi(CAMLine_11_io_wi),
    .io_key(CAMLine_11_io_key),
    .io_din(CAMLine_11_io_din),
    .io_hit(CAMLine_11_io_hit)
  );
  CAMLine CAMLine_12 ( // @[cam.scala 81:36]
    .clock(CAMLine_12_clock),
    .io_we(CAMLine_12_io_we),
    .io_wi(CAMLine_12_io_wi),
    .io_key(CAMLine_12_io_key),
    .io_din(CAMLine_12_io_din),
    .io_hit(CAMLine_12_io_hit)
  );
  CAMLine CAMLine_13 ( // @[cam.scala 81:36]
    .clock(CAMLine_13_clock),
    .io_we(CAMLine_13_io_we),
    .io_wi(CAMLine_13_io_wi),
    .io_key(CAMLine_13_io_key),
    .io_din(CAMLine_13_io_din),
    .io_hit(CAMLine_13_io_hit)
  );
  CAMLine CAMLine_14 ( // @[cam.scala 81:36]
    .clock(CAMLine_14_clock),
    .io_we(CAMLine_14_io_we),
    .io_wi(CAMLine_14_io_wi),
    .io_key(CAMLine_14_io_key),
    .io_din(CAMLine_14_io_din),
    .io_hit(CAMLine_14_io_hit)
  );
  CAMLine CAMLine_15 ( // @[cam.scala 81:36]
    .clock(CAMLine_15_clock),
    .io_we(CAMLine_15_io_we),
    .io_wi(CAMLine_15_io_wi),
    .io_key(CAMLine_15_io_key),
    .io_din(CAMLine_15_io_din),
    .io_hit(CAMLine_15_io_hit)
  );
  CAMLine CAMLine_16 ( // @[cam.scala 81:36]
    .clock(CAMLine_16_clock),
    .io_we(CAMLine_16_io_we),
    .io_wi(CAMLine_16_io_wi),
    .io_key(CAMLine_16_io_key),
    .io_din(CAMLine_16_io_din),
    .io_hit(CAMLine_16_io_hit)
  );
  CAMLine CAMLine_17 ( // @[cam.scala 81:36]
    .clock(CAMLine_17_clock),
    .io_we(CAMLine_17_io_we),
    .io_wi(CAMLine_17_io_wi),
    .io_key(CAMLine_17_io_key),
    .io_din(CAMLine_17_io_din),
    .io_hit(CAMLine_17_io_hit)
  );
  CAMLine CAMLine_18 ( // @[cam.scala 81:36]
    .clock(CAMLine_18_clock),
    .io_we(CAMLine_18_io_we),
    .io_wi(CAMLine_18_io_wi),
    .io_key(CAMLine_18_io_key),
    .io_din(CAMLine_18_io_din),
    .io_hit(CAMLine_18_io_hit)
  );
  CAMLine CAMLine_19 ( // @[cam.scala 81:36]
    .clock(CAMLine_19_clock),
    .io_we(CAMLine_19_io_we),
    .io_wi(CAMLine_19_io_wi),
    .io_key(CAMLine_19_io_key),
    .io_din(CAMLine_19_io_din),
    .io_hit(CAMLine_19_io_hit)
  );
  CAMLine CAMLine_20 ( // @[cam.scala 81:36]
    .clock(CAMLine_20_clock),
    .io_we(CAMLine_20_io_we),
    .io_wi(CAMLine_20_io_wi),
    .io_key(CAMLine_20_io_key),
    .io_din(CAMLine_20_io_din),
    .io_hit(CAMLine_20_io_hit)
  );
  CAMLine CAMLine_21 ( // @[cam.scala 81:36]
    .clock(CAMLine_21_clock),
    .io_we(CAMLine_21_io_we),
    .io_wi(CAMLine_21_io_wi),
    .io_key(CAMLine_21_io_key),
    .io_din(CAMLine_21_io_din),
    .io_hit(CAMLine_21_io_hit)
  );
  CAMLine CAMLine_22 ( // @[cam.scala 81:36]
    .clock(CAMLine_22_clock),
    .io_we(CAMLine_22_io_we),
    .io_wi(CAMLine_22_io_wi),
    .io_key(CAMLine_22_io_key),
    .io_din(CAMLine_22_io_din),
    .io_hit(CAMLine_22_io_hit)
  );
  CAMLine CAMLine_23 ( // @[cam.scala 81:36]
    .clock(CAMLine_23_clock),
    .io_we(CAMLine_23_io_we),
    .io_wi(CAMLine_23_io_wi),
    .io_key(CAMLine_23_io_key),
    .io_din(CAMLine_23_io_din),
    .io_hit(CAMLine_23_io_hit)
  );
  CAMLine CAMLine_24 ( // @[cam.scala 81:36]
    .clock(CAMLine_24_clock),
    .io_we(CAMLine_24_io_we),
    .io_wi(CAMLine_24_io_wi),
    .io_key(CAMLine_24_io_key),
    .io_din(CAMLine_24_io_din),
    .io_hit(CAMLine_24_io_hit)
  );
  CAMLine CAMLine_25 ( // @[cam.scala 81:36]
    .clock(CAMLine_25_clock),
    .io_we(CAMLine_25_io_we),
    .io_wi(CAMLine_25_io_wi),
    .io_key(CAMLine_25_io_key),
    .io_din(CAMLine_25_io_din),
    .io_hit(CAMLine_25_io_hit)
  );
  CAMLine CAMLine_26 ( // @[cam.scala 81:36]
    .clock(CAMLine_26_clock),
    .io_we(CAMLine_26_io_we),
    .io_wi(CAMLine_26_io_wi),
    .io_key(CAMLine_26_io_key),
    .io_din(CAMLine_26_io_din),
    .io_hit(CAMLine_26_io_hit)
  );
  CAMLine CAMLine_27 ( // @[cam.scala 81:36]
    .clock(CAMLine_27_clock),
    .io_we(CAMLine_27_io_we),
    .io_wi(CAMLine_27_io_wi),
    .io_key(CAMLine_27_io_key),
    .io_din(CAMLine_27_io_din),
    .io_hit(CAMLine_27_io_hit)
  );
  CAMLine CAMLine_28 ( // @[cam.scala 81:36]
    .clock(CAMLine_28_clock),
    .io_we(CAMLine_28_io_we),
    .io_wi(CAMLine_28_io_wi),
    .io_key(CAMLine_28_io_key),
    .io_din(CAMLine_28_io_din),
    .io_hit(CAMLine_28_io_hit)
  );
  CAMLine CAMLine_29 ( // @[cam.scala 81:36]
    .clock(CAMLine_29_clock),
    .io_we(CAMLine_29_io_we),
    .io_wi(CAMLine_29_io_wi),
    .io_key(CAMLine_29_io_key),
    .io_din(CAMLine_29_io_din),
    .io_hit(CAMLine_29_io_hit)
  );
  CAMLine CAMLine_30 ( // @[cam.scala 81:36]
    .clock(CAMLine_30_clock),
    .io_we(CAMLine_30_io_we),
    .io_wi(CAMLine_30_io_wi),
    .io_key(CAMLine_30_io_key),
    .io_din(CAMLine_30_io_din),
    .io_hit(CAMLine_30_io_hit)
  );
  CAMLine CAMLine_31 ( // @[cam.scala 81:36]
    .clock(CAMLine_31_clock),
    .io_we(CAMLine_31_io_we),
    .io_wi(CAMLine_31_io_wi),
    .io_key(CAMLine_31_io_key),
    .io_din(CAMLine_31_io_din),
    .io_hit(CAMLine_31_io_hit)
  );
  CAMLine CAMLine_32 ( // @[cam.scala 81:36]
    .clock(CAMLine_32_clock),
    .io_we(CAMLine_32_io_we),
    .io_wi(CAMLine_32_io_wi),
    .io_key(CAMLine_32_io_key),
    .io_din(CAMLine_32_io_din),
    .io_hit(CAMLine_32_io_hit)
  );
  CAMLine CAMLine_33 ( // @[cam.scala 81:36]
    .clock(CAMLine_33_clock),
    .io_we(CAMLine_33_io_we),
    .io_wi(CAMLine_33_io_wi),
    .io_key(CAMLine_33_io_key),
    .io_din(CAMLine_33_io_din),
    .io_hit(CAMLine_33_io_hit)
  );
  CAMLine CAMLine_34 ( // @[cam.scala 81:36]
    .clock(CAMLine_34_clock),
    .io_we(CAMLine_34_io_we),
    .io_wi(CAMLine_34_io_wi),
    .io_key(CAMLine_34_io_key),
    .io_din(CAMLine_34_io_din),
    .io_hit(CAMLine_34_io_hit)
  );
  CAMLine CAMLine_35 ( // @[cam.scala 81:36]
    .clock(CAMLine_35_clock),
    .io_we(CAMLine_35_io_we),
    .io_wi(CAMLine_35_io_wi),
    .io_key(CAMLine_35_io_key),
    .io_din(CAMLine_35_io_din),
    .io_hit(CAMLine_35_io_hit)
  );
  CAMLine CAMLine_36 ( // @[cam.scala 81:36]
    .clock(CAMLine_36_clock),
    .io_we(CAMLine_36_io_we),
    .io_wi(CAMLine_36_io_wi),
    .io_key(CAMLine_36_io_key),
    .io_din(CAMLine_36_io_din),
    .io_hit(CAMLine_36_io_hit)
  );
  CAMLine CAMLine_37 ( // @[cam.scala 81:36]
    .clock(CAMLine_37_clock),
    .io_we(CAMLine_37_io_we),
    .io_wi(CAMLine_37_io_wi),
    .io_key(CAMLine_37_io_key),
    .io_din(CAMLine_37_io_din),
    .io_hit(CAMLine_37_io_hit)
  );
  CAMLine CAMLine_38 ( // @[cam.scala 81:36]
    .clock(CAMLine_38_clock),
    .io_we(CAMLine_38_io_we),
    .io_wi(CAMLine_38_io_wi),
    .io_key(CAMLine_38_io_key),
    .io_din(CAMLine_38_io_din),
    .io_hit(CAMLine_38_io_hit)
  );
  CAMLine CAMLine_39 ( // @[cam.scala 81:36]
    .clock(CAMLine_39_clock),
    .io_we(CAMLine_39_io_we),
    .io_wi(CAMLine_39_io_wi),
    .io_key(CAMLine_39_io_key),
    .io_din(CAMLine_39_io_din),
    .io_hit(CAMLine_39_io_hit)
  );
  CAMLine CAMLine_40 ( // @[cam.scala 81:36]
    .clock(CAMLine_40_clock),
    .io_we(CAMLine_40_io_we),
    .io_wi(CAMLine_40_io_wi),
    .io_key(CAMLine_40_io_key),
    .io_din(CAMLine_40_io_din),
    .io_hit(CAMLine_40_io_hit)
  );
  CAMLine CAMLine_41 ( // @[cam.scala 81:36]
    .clock(CAMLine_41_clock),
    .io_we(CAMLine_41_io_we),
    .io_wi(CAMLine_41_io_wi),
    .io_key(CAMLine_41_io_key),
    .io_din(CAMLine_41_io_din),
    .io_hit(CAMLine_41_io_hit)
  );
  CAMLine CAMLine_42 ( // @[cam.scala 81:36]
    .clock(CAMLine_42_clock),
    .io_we(CAMLine_42_io_we),
    .io_wi(CAMLine_42_io_wi),
    .io_key(CAMLine_42_io_key),
    .io_din(CAMLine_42_io_din),
    .io_hit(CAMLine_42_io_hit)
  );
  CAMLine CAMLine_43 ( // @[cam.scala 81:36]
    .clock(CAMLine_43_clock),
    .io_we(CAMLine_43_io_we),
    .io_wi(CAMLine_43_io_wi),
    .io_key(CAMLine_43_io_key),
    .io_din(CAMLine_43_io_din),
    .io_hit(CAMLine_43_io_hit)
  );
  CAMLine CAMLine_44 ( // @[cam.scala 81:36]
    .clock(CAMLine_44_clock),
    .io_we(CAMLine_44_io_we),
    .io_wi(CAMLine_44_io_wi),
    .io_key(CAMLine_44_io_key),
    .io_din(CAMLine_44_io_din),
    .io_hit(CAMLine_44_io_hit)
  );
  CAMLine CAMLine_45 ( // @[cam.scala 81:36]
    .clock(CAMLine_45_clock),
    .io_we(CAMLine_45_io_we),
    .io_wi(CAMLine_45_io_wi),
    .io_key(CAMLine_45_io_key),
    .io_din(CAMLine_45_io_din),
    .io_hit(CAMLine_45_io_hit)
  );
  CAMLine CAMLine_46 ( // @[cam.scala 81:36]
    .clock(CAMLine_46_clock),
    .io_we(CAMLine_46_io_we),
    .io_wi(CAMLine_46_io_wi),
    .io_key(CAMLine_46_io_key),
    .io_din(CAMLine_46_io_din),
    .io_hit(CAMLine_46_io_hit)
  );
  CAMLine CAMLine_47 ( // @[cam.scala 81:36]
    .clock(CAMLine_47_clock),
    .io_we(CAMLine_47_io_we),
    .io_wi(CAMLine_47_io_wi),
    .io_key(CAMLine_47_io_key),
    .io_din(CAMLine_47_io_din),
    .io_hit(CAMLine_47_io_hit)
  );
  CAMLine CAMLine_48 ( // @[cam.scala 81:36]
    .clock(CAMLine_48_clock),
    .io_we(CAMLine_48_io_we),
    .io_wi(CAMLine_48_io_wi),
    .io_key(CAMLine_48_io_key),
    .io_din(CAMLine_48_io_din),
    .io_hit(CAMLine_48_io_hit)
  );
  CAMLine CAMLine_49 ( // @[cam.scala 81:36]
    .clock(CAMLine_49_clock),
    .io_we(CAMLine_49_io_we),
    .io_wi(CAMLine_49_io_wi),
    .io_key(CAMLine_49_io_key),
    .io_din(CAMLine_49_io_din),
    .io_hit(CAMLine_49_io_hit)
  );
  CAMLine CAMLine_50 ( // @[cam.scala 81:36]
    .clock(CAMLine_50_clock),
    .io_we(CAMLine_50_io_we),
    .io_wi(CAMLine_50_io_wi),
    .io_key(CAMLine_50_io_key),
    .io_din(CAMLine_50_io_din),
    .io_hit(CAMLine_50_io_hit)
  );
  CAMLine CAMLine_51 ( // @[cam.scala 81:36]
    .clock(CAMLine_51_clock),
    .io_we(CAMLine_51_io_we),
    .io_wi(CAMLine_51_io_wi),
    .io_key(CAMLine_51_io_key),
    .io_din(CAMLine_51_io_din),
    .io_hit(CAMLine_51_io_hit)
  );
  CAMLine CAMLine_52 ( // @[cam.scala 81:36]
    .clock(CAMLine_52_clock),
    .io_we(CAMLine_52_io_we),
    .io_wi(CAMLine_52_io_wi),
    .io_key(CAMLine_52_io_key),
    .io_din(CAMLine_52_io_din),
    .io_hit(CAMLine_52_io_hit)
  );
  CAMLine CAMLine_53 ( // @[cam.scala 81:36]
    .clock(CAMLine_53_clock),
    .io_we(CAMLine_53_io_we),
    .io_wi(CAMLine_53_io_wi),
    .io_key(CAMLine_53_io_key),
    .io_din(CAMLine_53_io_din),
    .io_hit(CAMLine_53_io_hit)
  );
  CAMLine CAMLine_54 ( // @[cam.scala 81:36]
    .clock(CAMLine_54_clock),
    .io_we(CAMLine_54_io_we),
    .io_wi(CAMLine_54_io_wi),
    .io_key(CAMLine_54_io_key),
    .io_din(CAMLine_54_io_din),
    .io_hit(CAMLine_54_io_hit)
  );
  CAMLine CAMLine_55 ( // @[cam.scala 81:36]
    .clock(CAMLine_55_clock),
    .io_we(CAMLine_55_io_we),
    .io_wi(CAMLine_55_io_wi),
    .io_key(CAMLine_55_io_key),
    .io_din(CAMLine_55_io_din),
    .io_hit(CAMLine_55_io_hit)
  );
  CAMLine CAMLine_56 ( // @[cam.scala 81:36]
    .clock(CAMLine_56_clock),
    .io_we(CAMLine_56_io_we),
    .io_wi(CAMLine_56_io_wi),
    .io_key(CAMLine_56_io_key),
    .io_din(CAMLine_56_io_din),
    .io_hit(CAMLine_56_io_hit)
  );
  CAMLine CAMLine_57 ( // @[cam.scala 81:36]
    .clock(CAMLine_57_clock),
    .io_we(CAMLine_57_io_we),
    .io_wi(CAMLine_57_io_wi),
    .io_key(CAMLine_57_io_key),
    .io_din(CAMLine_57_io_din),
    .io_hit(CAMLine_57_io_hit)
  );
  CAMLine CAMLine_58 ( // @[cam.scala 81:36]
    .clock(CAMLine_58_clock),
    .io_we(CAMLine_58_io_we),
    .io_wi(CAMLine_58_io_wi),
    .io_key(CAMLine_58_io_key),
    .io_din(CAMLine_58_io_din),
    .io_hit(CAMLine_58_io_hit)
  );
  CAMLine CAMLine_59 ( // @[cam.scala 81:36]
    .clock(CAMLine_59_clock),
    .io_we(CAMLine_59_io_we),
    .io_wi(CAMLine_59_io_wi),
    .io_key(CAMLine_59_io_key),
    .io_din(CAMLine_59_io_din),
    .io_hit(CAMLine_59_io_hit)
  );
  CAMLine CAMLine_60 ( // @[cam.scala 81:36]
    .clock(CAMLine_60_clock),
    .io_we(CAMLine_60_io_we),
    .io_wi(CAMLine_60_io_wi),
    .io_key(CAMLine_60_io_key),
    .io_din(CAMLine_60_io_din),
    .io_hit(CAMLine_60_io_hit)
  );
  CAMLine CAMLine_61 ( // @[cam.scala 81:36]
    .clock(CAMLine_61_clock),
    .io_we(CAMLine_61_io_we),
    .io_wi(CAMLine_61_io_wi),
    .io_key(CAMLine_61_io_key),
    .io_din(CAMLine_61_io_din),
    .io_hit(CAMLine_61_io_hit)
  );
  CAMLine CAMLine_62 ( // @[cam.scala 81:36]
    .clock(CAMLine_62_clock),
    .io_we(CAMLine_62_io_we),
    .io_wi(CAMLine_62_io_wi),
    .io_key(CAMLine_62_io_key),
    .io_din(CAMLine_62_io_din),
    .io_hit(CAMLine_62_io_hit)
  );
  CAMLine CAMLine_63 ( // @[cam.scala 81:36]
    .clock(CAMLine_63_clock),
    .io_we(CAMLine_63_io_we),
    .io_wi(CAMLine_63_io_wi),
    .io_key(CAMLine_63_io_key),
    .io_din(CAMLine_63_io_din),
    .io_hit(CAMLine_63_io_hit)
  );
  CAMLine CAMLine_64 ( // @[cam.scala 81:36]
    .clock(CAMLine_64_clock),
    .io_we(CAMLine_64_io_we),
    .io_wi(CAMLine_64_io_wi),
    .io_key(CAMLine_64_io_key),
    .io_din(CAMLine_64_io_din),
    .io_hit(CAMLine_64_io_hit)
  );
  CAMLine CAMLine_65 ( // @[cam.scala 81:36]
    .clock(CAMLine_65_clock),
    .io_we(CAMLine_65_io_we),
    .io_wi(CAMLine_65_io_wi),
    .io_key(CAMLine_65_io_key),
    .io_din(CAMLine_65_io_din),
    .io_hit(CAMLine_65_io_hit)
  );
  CAMLine CAMLine_66 ( // @[cam.scala 81:36]
    .clock(CAMLine_66_clock),
    .io_we(CAMLine_66_io_we),
    .io_wi(CAMLine_66_io_wi),
    .io_key(CAMLine_66_io_key),
    .io_din(CAMLine_66_io_din),
    .io_hit(CAMLine_66_io_hit)
  );
  CAMLine CAMLine_67 ( // @[cam.scala 81:36]
    .clock(CAMLine_67_clock),
    .io_we(CAMLine_67_io_we),
    .io_wi(CAMLine_67_io_wi),
    .io_key(CAMLine_67_io_key),
    .io_din(CAMLine_67_io_din),
    .io_hit(CAMLine_67_io_hit)
  );
  CAMLine CAMLine_68 ( // @[cam.scala 81:36]
    .clock(CAMLine_68_clock),
    .io_we(CAMLine_68_io_we),
    .io_wi(CAMLine_68_io_wi),
    .io_key(CAMLine_68_io_key),
    .io_din(CAMLine_68_io_din),
    .io_hit(CAMLine_68_io_hit)
  );
  CAMLine CAMLine_69 ( // @[cam.scala 81:36]
    .clock(CAMLine_69_clock),
    .io_we(CAMLine_69_io_we),
    .io_wi(CAMLine_69_io_wi),
    .io_key(CAMLine_69_io_key),
    .io_din(CAMLine_69_io_din),
    .io_hit(CAMLine_69_io_hit)
  );
  CAMLine CAMLine_70 ( // @[cam.scala 81:36]
    .clock(CAMLine_70_clock),
    .io_we(CAMLine_70_io_we),
    .io_wi(CAMLine_70_io_wi),
    .io_key(CAMLine_70_io_key),
    .io_din(CAMLine_70_io_din),
    .io_hit(CAMLine_70_io_hit)
  );
  CAMLine CAMLine_71 ( // @[cam.scala 81:36]
    .clock(CAMLine_71_clock),
    .io_we(CAMLine_71_io_we),
    .io_wi(CAMLine_71_io_wi),
    .io_key(CAMLine_71_io_key),
    .io_din(CAMLine_71_io_din),
    .io_hit(CAMLine_71_io_hit)
  );
  CAMLine CAMLine_72 ( // @[cam.scala 81:36]
    .clock(CAMLine_72_clock),
    .io_we(CAMLine_72_io_we),
    .io_wi(CAMLine_72_io_wi),
    .io_key(CAMLine_72_io_key),
    .io_din(CAMLine_72_io_din),
    .io_hit(CAMLine_72_io_hit)
  );
  CAMLine CAMLine_73 ( // @[cam.scala 81:36]
    .clock(CAMLine_73_clock),
    .io_we(CAMLine_73_io_we),
    .io_wi(CAMLine_73_io_wi),
    .io_key(CAMLine_73_io_key),
    .io_din(CAMLine_73_io_din),
    .io_hit(CAMLine_73_io_hit)
  );
  CAMLine CAMLine_74 ( // @[cam.scala 81:36]
    .clock(CAMLine_74_clock),
    .io_we(CAMLine_74_io_we),
    .io_wi(CAMLine_74_io_wi),
    .io_key(CAMLine_74_io_key),
    .io_din(CAMLine_74_io_din),
    .io_hit(CAMLine_74_io_hit)
  );
  CAMLine CAMLine_75 ( // @[cam.scala 81:36]
    .clock(CAMLine_75_clock),
    .io_we(CAMLine_75_io_we),
    .io_wi(CAMLine_75_io_wi),
    .io_key(CAMLine_75_io_key),
    .io_din(CAMLine_75_io_din),
    .io_hit(CAMLine_75_io_hit)
  );
  CAMLine CAMLine_76 ( // @[cam.scala 81:36]
    .clock(CAMLine_76_clock),
    .io_we(CAMLine_76_io_we),
    .io_wi(CAMLine_76_io_wi),
    .io_key(CAMLine_76_io_key),
    .io_din(CAMLine_76_io_din),
    .io_hit(CAMLine_76_io_hit)
  );
  CAMLine CAMLine_77 ( // @[cam.scala 81:36]
    .clock(CAMLine_77_clock),
    .io_we(CAMLine_77_io_we),
    .io_wi(CAMLine_77_io_wi),
    .io_key(CAMLine_77_io_key),
    .io_din(CAMLine_77_io_din),
    .io_hit(CAMLine_77_io_hit)
  );
  CAMLine CAMLine_78 ( // @[cam.scala 81:36]
    .clock(CAMLine_78_clock),
    .io_we(CAMLine_78_io_we),
    .io_wi(CAMLine_78_io_wi),
    .io_key(CAMLine_78_io_key),
    .io_din(CAMLine_78_io_din),
    .io_hit(CAMLine_78_io_hit)
  );
  CAMLine CAMLine_79 ( // @[cam.scala 81:36]
    .clock(CAMLine_79_clock),
    .io_we(CAMLine_79_io_we),
    .io_wi(CAMLine_79_io_wi),
    .io_key(CAMLine_79_io_key),
    .io_din(CAMLine_79_io_din),
    .io_hit(CAMLine_79_io_hit)
  );
  CAMLine CAMLine_80 ( // @[cam.scala 81:36]
    .clock(CAMLine_80_clock),
    .io_we(CAMLine_80_io_we),
    .io_wi(CAMLine_80_io_wi),
    .io_key(CAMLine_80_io_key),
    .io_din(CAMLine_80_io_din),
    .io_hit(CAMLine_80_io_hit)
  );
  CAMLine CAMLine_81 ( // @[cam.scala 81:36]
    .clock(CAMLine_81_clock),
    .io_we(CAMLine_81_io_we),
    .io_wi(CAMLine_81_io_wi),
    .io_key(CAMLine_81_io_key),
    .io_din(CAMLine_81_io_din),
    .io_hit(CAMLine_81_io_hit)
  );
  CAMLine CAMLine_82 ( // @[cam.scala 81:36]
    .clock(CAMLine_82_clock),
    .io_we(CAMLine_82_io_we),
    .io_wi(CAMLine_82_io_wi),
    .io_key(CAMLine_82_io_key),
    .io_din(CAMLine_82_io_din),
    .io_hit(CAMLine_82_io_hit)
  );
  CAMLine CAMLine_83 ( // @[cam.scala 81:36]
    .clock(CAMLine_83_clock),
    .io_we(CAMLine_83_io_we),
    .io_wi(CAMLine_83_io_wi),
    .io_key(CAMLine_83_io_key),
    .io_din(CAMLine_83_io_din),
    .io_hit(CAMLine_83_io_hit)
  );
  CAMLine CAMLine_84 ( // @[cam.scala 81:36]
    .clock(CAMLine_84_clock),
    .io_we(CAMLine_84_io_we),
    .io_wi(CAMLine_84_io_wi),
    .io_key(CAMLine_84_io_key),
    .io_din(CAMLine_84_io_din),
    .io_hit(CAMLine_84_io_hit)
  );
  CAMLine CAMLine_85 ( // @[cam.scala 81:36]
    .clock(CAMLine_85_clock),
    .io_we(CAMLine_85_io_we),
    .io_wi(CAMLine_85_io_wi),
    .io_key(CAMLine_85_io_key),
    .io_din(CAMLine_85_io_din),
    .io_hit(CAMLine_85_io_hit)
  );
  CAMLine CAMLine_86 ( // @[cam.scala 81:36]
    .clock(CAMLine_86_clock),
    .io_we(CAMLine_86_io_we),
    .io_wi(CAMLine_86_io_wi),
    .io_key(CAMLine_86_io_key),
    .io_din(CAMLine_86_io_din),
    .io_hit(CAMLine_86_io_hit)
  );
  CAMLine CAMLine_87 ( // @[cam.scala 81:36]
    .clock(CAMLine_87_clock),
    .io_we(CAMLine_87_io_we),
    .io_wi(CAMLine_87_io_wi),
    .io_key(CAMLine_87_io_key),
    .io_din(CAMLine_87_io_din),
    .io_hit(CAMLine_87_io_hit)
  );
  CAMLine CAMLine_88 ( // @[cam.scala 81:36]
    .clock(CAMLine_88_clock),
    .io_we(CAMLine_88_io_we),
    .io_wi(CAMLine_88_io_wi),
    .io_key(CAMLine_88_io_key),
    .io_din(CAMLine_88_io_din),
    .io_hit(CAMLine_88_io_hit)
  );
  CAMLine CAMLine_89 ( // @[cam.scala 81:36]
    .clock(CAMLine_89_clock),
    .io_we(CAMLine_89_io_we),
    .io_wi(CAMLine_89_io_wi),
    .io_key(CAMLine_89_io_key),
    .io_din(CAMLine_89_io_din),
    .io_hit(CAMLine_89_io_hit)
  );
  CAMLine CAMLine_90 ( // @[cam.scala 81:36]
    .clock(CAMLine_90_clock),
    .io_we(CAMLine_90_io_we),
    .io_wi(CAMLine_90_io_wi),
    .io_key(CAMLine_90_io_key),
    .io_din(CAMLine_90_io_din),
    .io_hit(CAMLine_90_io_hit)
  );
  CAMLine CAMLine_91 ( // @[cam.scala 81:36]
    .clock(CAMLine_91_clock),
    .io_we(CAMLine_91_io_we),
    .io_wi(CAMLine_91_io_wi),
    .io_key(CAMLine_91_io_key),
    .io_din(CAMLine_91_io_din),
    .io_hit(CAMLine_91_io_hit)
  );
  CAMLine CAMLine_92 ( // @[cam.scala 81:36]
    .clock(CAMLine_92_clock),
    .io_we(CAMLine_92_io_we),
    .io_wi(CAMLine_92_io_wi),
    .io_key(CAMLine_92_io_key),
    .io_din(CAMLine_92_io_din),
    .io_hit(CAMLine_92_io_hit)
  );
  CAMLine CAMLine_93 ( // @[cam.scala 81:36]
    .clock(CAMLine_93_clock),
    .io_we(CAMLine_93_io_we),
    .io_wi(CAMLine_93_io_wi),
    .io_key(CAMLine_93_io_key),
    .io_din(CAMLine_93_io_din),
    .io_hit(CAMLine_93_io_hit)
  );
  CAMLine CAMLine_94 ( // @[cam.scala 81:36]
    .clock(CAMLine_94_clock),
    .io_we(CAMLine_94_io_we),
    .io_wi(CAMLine_94_io_wi),
    .io_key(CAMLine_94_io_key),
    .io_din(CAMLine_94_io_din),
    .io_hit(CAMLine_94_io_hit)
  );
  CAMLine CAMLine_95 ( // @[cam.scala 81:36]
    .clock(CAMLine_95_clock),
    .io_we(CAMLine_95_io_we),
    .io_wi(CAMLine_95_io_wi),
    .io_key(CAMLine_95_io_key),
    .io_din(CAMLine_95_io_din),
    .io_hit(CAMLine_95_io_hit)
  );
  CAMLine CAMLine_96 ( // @[cam.scala 81:36]
    .clock(CAMLine_96_clock),
    .io_we(CAMLine_96_io_we),
    .io_wi(CAMLine_96_io_wi),
    .io_key(CAMLine_96_io_key),
    .io_din(CAMLine_96_io_din),
    .io_hit(CAMLine_96_io_hit)
  );
  CAMLine CAMLine_97 ( // @[cam.scala 81:36]
    .clock(CAMLine_97_clock),
    .io_we(CAMLine_97_io_we),
    .io_wi(CAMLine_97_io_wi),
    .io_key(CAMLine_97_io_key),
    .io_din(CAMLine_97_io_din),
    .io_hit(CAMLine_97_io_hit)
  );
  CAMLine CAMLine_98 ( // @[cam.scala 81:36]
    .clock(CAMLine_98_clock),
    .io_we(CAMLine_98_io_we),
    .io_wi(CAMLine_98_io_wi),
    .io_key(CAMLine_98_io_key),
    .io_din(CAMLine_98_io_din),
    .io_hit(CAMLine_98_io_hit)
  );
  CAMLine CAMLine_99 ( // @[cam.scala 81:36]
    .clock(CAMLine_99_clock),
    .io_we(CAMLine_99_io_we),
    .io_wi(CAMLine_99_io_wi),
    .io_key(CAMLine_99_io_key),
    .io_din(CAMLine_99_io_din),
    .io_hit(CAMLine_99_io_hit)
  );
  CAMLine CAMLine_100 ( // @[cam.scala 81:36]
    .clock(CAMLine_100_clock),
    .io_we(CAMLine_100_io_we),
    .io_wi(CAMLine_100_io_wi),
    .io_key(CAMLine_100_io_key),
    .io_din(CAMLine_100_io_din),
    .io_hit(CAMLine_100_io_hit)
  );
  CAMLine CAMLine_101 ( // @[cam.scala 81:36]
    .clock(CAMLine_101_clock),
    .io_we(CAMLine_101_io_we),
    .io_wi(CAMLine_101_io_wi),
    .io_key(CAMLine_101_io_key),
    .io_din(CAMLine_101_io_din),
    .io_hit(CAMLine_101_io_hit)
  );
  CAMLine CAMLine_102 ( // @[cam.scala 81:36]
    .clock(CAMLine_102_clock),
    .io_we(CAMLine_102_io_we),
    .io_wi(CAMLine_102_io_wi),
    .io_key(CAMLine_102_io_key),
    .io_din(CAMLine_102_io_din),
    .io_hit(CAMLine_102_io_hit)
  );
  CAMLine CAMLine_103 ( // @[cam.scala 81:36]
    .clock(CAMLine_103_clock),
    .io_we(CAMLine_103_io_we),
    .io_wi(CAMLine_103_io_wi),
    .io_key(CAMLine_103_io_key),
    .io_din(CAMLine_103_io_din),
    .io_hit(CAMLine_103_io_hit)
  );
  CAMLine CAMLine_104 ( // @[cam.scala 81:36]
    .clock(CAMLine_104_clock),
    .io_we(CAMLine_104_io_we),
    .io_wi(CAMLine_104_io_wi),
    .io_key(CAMLine_104_io_key),
    .io_din(CAMLine_104_io_din),
    .io_hit(CAMLine_104_io_hit)
  );
  CAMLine CAMLine_105 ( // @[cam.scala 81:36]
    .clock(CAMLine_105_clock),
    .io_we(CAMLine_105_io_we),
    .io_wi(CAMLine_105_io_wi),
    .io_key(CAMLine_105_io_key),
    .io_din(CAMLine_105_io_din),
    .io_hit(CAMLine_105_io_hit)
  );
  CAMLine CAMLine_106 ( // @[cam.scala 81:36]
    .clock(CAMLine_106_clock),
    .io_we(CAMLine_106_io_we),
    .io_wi(CAMLine_106_io_wi),
    .io_key(CAMLine_106_io_key),
    .io_din(CAMLine_106_io_din),
    .io_hit(CAMLine_106_io_hit)
  );
  CAMLine CAMLine_107 ( // @[cam.scala 81:36]
    .clock(CAMLine_107_clock),
    .io_we(CAMLine_107_io_we),
    .io_wi(CAMLine_107_io_wi),
    .io_key(CAMLine_107_io_key),
    .io_din(CAMLine_107_io_din),
    .io_hit(CAMLine_107_io_hit)
  );
  CAMLine CAMLine_108 ( // @[cam.scala 81:36]
    .clock(CAMLine_108_clock),
    .io_we(CAMLine_108_io_we),
    .io_wi(CAMLine_108_io_wi),
    .io_key(CAMLine_108_io_key),
    .io_din(CAMLine_108_io_din),
    .io_hit(CAMLine_108_io_hit)
  );
  CAMLine CAMLine_109 ( // @[cam.scala 81:36]
    .clock(CAMLine_109_clock),
    .io_we(CAMLine_109_io_we),
    .io_wi(CAMLine_109_io_wi),
    .io_key(CAMLine_109_io_key),
    .io_din(CAMLine_109_io_din),
    .io_hit(CAMLine_109_io_hit)
  );
  CAMLine CAMLine_110 ( // @[cam.scala 81:36]
    .clock(CAMLine_110_clock),
    .io_we(CAMLine_110_io_we),
    .io_wi(CAMLine_110_io_wi),
    .io_key(CAMLine_110_io_key),
    .io_din(CAMLine_110_io_din),
    .io_hit(CAMLine_110_io_hit)
  );
  CAMLine CAMLine_111 ( // @[cam.scala 81:36]
    .clock(CAMLine_111_clock),
    .io_we(CAMLine_111_io_we),
    .io_wi(CAMLine_111_io_wi),
    .io_key(CAMLine_111_io_key),
    .io_din(CAMLine_111_io_din),
    .io_hit(CAMLine_111_io_hit)
  );
  CAMLine CAMLine_112 ( // @[cam.scala 81:36]
    .clock(CAMLine_112_clock),
    .io_we(CAMLine_112_io_we),
    .io_wi(CAMLine_112_io_wi),
    .io_key(CAMLine_112_io_key),
    .io_din(CAMLine_112_io_din),
    .io_hit(CAMLine_112_io_hit)
  );
  CAMLine CAMLine_113 ( // @[cam.scala 81:36]
    .clock(CAMLine_113_clock),
    .io_we(CAMLine_113_io_we),
    .io_wi(CAMLine_113_io_wi),
    .io_key(CAMLine_113_io_key),
    .io_din(CAMLine_113_io_din),
    .io_hit(CAMLine_113_io_hit)
  );
  CAMLine CAMLine_114 ( // @[cam.scala 81:36]
    .clock(CAMLine_114_clock),
    .io_we(CAMLine_114_io_we),
    .io_wi(CAMLine_114_io_wi),
    .io_key(CAMLine_114_io_key),
    .io_din(CAMLine_114_io_din),
    .io_hit(CAMLine_114_io_hit)
  );
  CAMLine CAMLine_115 ( // @[cam.scala 81:36]
    .clock(CAMLine_115_clock),
    .io_we(CAMLine_115_io_we),
    .io_wi(CAMLine_115_io_wi),
    .io_key(CAMLine_115_io_key),
    .io_din(CAMLine_115_io_din),
    .io_hit(CAMLine_115_io_hit)
  );
  CAMLine CAMLine_116 ( // @[cam.scala 81:36]
    .clock(CAMLine_116_clock),
    .io_we(CAMLine_116_io_we),
    .io_wi(CAMLine_116_io_wi),
    .io_key(CAMLine_116_io_key),
    .io_din(CAMLine_116_io_din),
    .io_hit(CAMLine_116_io_hit)
  );
  CAMLine CAMLine_117 ( // @[cam.scala 81:36]
    .clock(CAMLine_117_clock),
    .io_we(CAMLine_117_io_we),
    .io_wi(CAMLine_117_io_wi),
    .io_key(CAMLine_117_io_key),
    .io_din(CAMLine_117_io_din),
    .io_hit(CAMLine_117_io_hit)
  );
  CAMLine CAMLine_118 ( // @[cam.scala 81:36]
    .clock(CAMLine_118_clock),
    .io_we(CAMLine_118_io_we),
    .io_wi(CAMLine_118_io_wi),
    .io_key(CAMLine_118_io_key),
    .io_din(CAMLine_118_io_din),
    .io_hit(CAMLine_118_io_hit)
  );
  CAMLine CAMLine_119 ( // @[cam.scala 81:36]
    .clock(CAMLine_119_clock),
    .io_we(CAMLine_119_io_we),
    .io_wi(CAMLine_119_io_wi),
    .io_key(CAMLine_119_io_key),
    .io_din(CAMLine_119_io_din),
    .io_hit(CAMLine_119_io_hit)
  );
  CAMLine CAMLine_120 ( // @[cam.scala 81:36]
    .clock(CAMLine_120_clock),
    .io_we(CAMLine_120_io_we),
    .io_wi(CAMLine_120_io_wi),
    .io_key(CAMLine_120_io_key),
    .io_din(CAMLine_120_io_din),
    .io_hit(CAMLine_120_io_hit)
  );
  CAMLine CAMLine_121 ( // @[cam.scala 81:36]
    .clock(CAMLine_121_clock),
    .io_we(CAMLine_121_io_we),
    .io_wi(CAMLine_121_io_wi),
    .io_key(CAMLine_121_io_key),
    .io_din(CAMLine_121_io_din),
    .io_hit(CAMLine_121_io_hit)
  );
  CAMLine CAMLine_122 ( // @[cam.scala 81:36]
    .clock(CAMLine_122_clock),
    .io_we(CAMLine_122_io_we),
    .io_wi(CAMLine_122_io_wi),
    .io_key(CAMLine_122_io_key),
    .io_din(CAMLine_122_io_din),
    .io_hit(CAMLine_122_io_hit)
  );
  CAMLine CAMLine_123 ( // @[cam.scala 81:36]
    .clock(CAMLine_123_clock),
    .io_we(CAMLine_123_io_we),
    .io_wi(CAMLine_123_io_wi),
    .io_key(CAMLine_123_io_key),
    .io_din(CAMLine_123_io_din),
    .io_hit(CAMLine_123_io_hit)
  );
  CAMLine CAMLine_124 ( // @[cam.scala 81:36]
    .clock(CAMLine_124_clock),
    .io_we(CAMLine_124_io_we),
    .io_wi(CAMLine_124_io_wi),
    .io_key(CAMLine_124_io_key),
    .io_din(CAMLine_124_io_din),
    .io_hit(CAMLine_124_io_hit)
  );
  CAMLine CAMLine_125 ( // @[cam.scala 81:36]
    .clock(CAMLine_125_clock),
    .io_we(CAMLine_125_io_we),
    .io_wi(CAMLine_125_io_wi),
    .io_key(CAMLine_125_io_key),
    .io_din(CAMLine_125_io_din),
    .io_hit(CAMLine_125_io_hit)
  );
  CAMLine CAMLine_126 ( // @[cam.scala 81:36]
    .clock(CAMLine_126_clock),
    .io_we(CAMLine_126_io_we),
    .io_wi(CAMLine_126_io_wi),
    .io_key(CAMLine_126_io_key),
    .io_din(CAMLine_126_io_din),
    .io_hit(CAMLine_126_io_hit)
  );
  CAMLine CAMLine_127 ( // @[cam.scala 81:36]
    .clock(CAMLine_127_clock),
    .io_we(CAMLine_127_io_we),
    .io_wi(CAMLine_127_io_wi),
    .io_key(CAMLine_127_io_key),
    .io_din(CAMLine_127_io_din),
    .io_hit(CAMLine_127_io_hit)
  );
  assign io_hit = _io_hit_T_119 | CAMLine_121_io_hit | CAMLine_122_io_hit | CAMLine_123_io_hit | CAMLine_124_io_hit |
    CAMLine_125_io_hit | CAMLine_126_io_hit | CAMLine_127_io_hit; // @[cam.scala 93:27]
  assign CAMLine_clock = clock;
  assign CAMLine_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_io_wi = io_waddr[0]; // @[cam.scala 86:31]
  assign CAMLine_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_1_clock = clock;
  assign CAMLine_1_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_1_io_wi = io_waddr[1]; // @[cam.scala 86:31]
  assign CAMLine_1_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_1_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_2_clock = clock;
  assign CAMLine_2_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_2_io_wi = io_waddr[2]; // @[cam.scala 86:31]
  assign CAMLine_2_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_2_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_3_clock = clock;
  assign CAMLine_3_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_3_io_wi = io_waddr[3]; // @[cam.scala 86:31]
  assign CAMLine_3_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_3_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_4_clock = clock;
  assign CAMLine_4_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_4_io_wi = io_waddr[4]; // @[cam.scala 86:31]
  assign CAMLine_4_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_4_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_5_clock = clock;
  assign CAMLine_5_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_5_io_wi = io_waddr[5]; // @[cam.scala 86:31]
  assign CAMLine_5_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_5_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_6_clock = clock;
  assign CAMLine_6_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_6_io_wi = io_waddr[6]; // @[cam.scala 86:31]
  assign CAMLine_6_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_6_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_7_clock = clock;
  assign CAMLine_7_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_7_io_wi = io_waddr[7]; // @[cam.scala 86:31]
  assign CAMLine_7_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_7_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_8_clock = clock;
  assign CAMLine_8_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_8_io_wi = io_waddr[8]; // @[cam.scala 86:31]
  assign CAMLine_8_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_8_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_9_clock = clock;
  assign CAMLine_9_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_9_io_wi = io_waddr[9]; // @[cam.scala 86:31]
  assign CAMLine_9_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_9_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_10_clock = clock;
  assign CAMLine_10_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_10_io_wi = io_waddr[10]; // @[cam.scala 86:31]
  assign CAMLine_10_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_10_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_11_clock = clock;
  assign CAMLine_11_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_11_io_wi = io_waddr[11]; // @[cam.scala 86:31]
  assign CAMLine_11_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_11_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_12_clock = clock;
  assign CAMLine_12_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_12_io_wi = io_waddr[12]; // @[cam.scala 86:31]
  assign CAMLine_12_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_12_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_13_clock = clock;
  assign CAMLine_13_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_13_io_wi = io_waddr[13]; // @[cam.scala 86:31]
  assign CAMLine_13_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_13_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_14_clock = clock;
  assign CAMLine_14_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_14_io_wi = io_waddr[14]; // @[cam.scala 86:31]
  assign CAMLine_14_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_14_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_15_clock = clock;
  assign CAMLine_15_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_15_io_wi = io_waddr[15]; // @[cam.scala 86:31]
  assign CAMLine_15_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_15_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_16_clock = clock;
  assign CAMLine_16_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_16_io_wi = io_waddr[16]; // @[cam.scala 86:31]
  assign CAMLine_16_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_16_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_17_clock = clock;
  assign CAMLine_17_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_17_io_wi = io_waddr[17]; // @[cam.scala 86:31]
  assign CAMLine_17_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_17_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_18_clock = clock;
  assign CAMLine_18_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_18_io_wi = io_waddr[18]; // @[cam.scala 86:31]
  assign CAMLine_18_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_18_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_19_clock = clock;
  assign CAMLine_19_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_19_io_wi = io_waddr[19]; // @[cam.scala 86:31]
  assign CAMLine_19_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_19_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_20_clock = clock;
  assign CAMLine_20_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_20_io_wi = io_waddr[20]; // @[cam.scala 86:31]
  assign CAMLine_20_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_20_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_21_clock = clock;
  assign CAMLine_21_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_21_io_wi = io_waddr[21]; // @[cam.scala 86:31]
  assign CAMLine_21_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_21_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_22_clock = clock;
  assign CAMLine_22_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_22_io_wi = io_waddr[22]; // @[cam.scala 86:31]
  assign CAMLine_22_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_22_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_23_clock = clock;
  assign CAMLine_23_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_23_io_wi = io_waddr[23]; // @[cam.scala 86:31]
  assign CAMLine_23_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_23_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_24_clock = clock;
  assign CAMLine_24_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_24_io_wi = io_waddr[24]; // @[cam.scala 86:31]
  assign CAMLine_24_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_24_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_25_clock = clock;
  assign CAMLine_25_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_25_io_wi = io_waddr[25]; // @[cam.scala 86:31]
  assign CAMLine_25_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_25_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_26_clock = clock;
  assign CAMLine_26_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_26_io_wi = io_waddr[26]; // @[cam.scala 86:31]
  assign CAMLine_26_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_26_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_27_clock = clock;
  assign CAMLine_27_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_27_io_wi = io_waddr[27]; // @[cam.scala 86:31]
  assign CAMLine_27_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_27_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_28_clock = clock;
  assign CAMLine_28_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_28_io_wi = io_waddr[28]; // @[cam.scala 86:31]
  assign CAMLine_28_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_28_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_29_clock = clock;
  assign CAMLine_29_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_29_io_wi = io_waddr[29]; // @[cam.scala 86:31]
  assign CAMLine_29_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_29_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_30_clock = clock;
  assign CAMLine_30_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_30_io_wi = io_waddr[30]; // @[cam.scala 86:31]
  assign CAMLine_30_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_30_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_31_clock = clock;
  assign CAMLine_31_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_31_io_wi = io_waddr[31]; // @[cam.scala 86:31]
  assign CAMLine_31_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_31_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_32_clock = clock;
  assign CAMLine_32_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_32_io_wi = io_waddr[32]; // @[cam.scala 86:31]
  assign CAMLine_32_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_32_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_33_clock = clock;
  assign CAMLine_33_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_33_io_wi = io_waddr[33]; // @[cam.scala 86:31]
  assign CAMLine_33_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_33_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_34_clock = clock;
  assign CAMLine_34_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_34_io_wi = io_waddr[34]; // @[cam.scala 86:31]
  assign CAMLine_34_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_34_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_35_clock = clock;
  assign CAMLine_35_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_35_io_wi = io_waddr[35]; // @[cam.scala 86:31]
  assign CAMLine_35_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_35_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_36_clock = clock;
  assign CAMLine_36_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_36_io_wi = io_waddr[36]; // @[cam.scala 86:31]
  assign CAMLine_36_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_36_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_37_clock = clock;
  assign CAMLine_37_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_37_io_wi = io_waddr[37]; // @[cam.scala 86:31]
  assign CAMLine_37_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_37_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_38_clock = clock;
  assign CAMLine_38_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_38_io_wi = io_waddr[38]; // @[cam.scala 86:31]
  assign CAMLine_38_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_38_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_39_clock = clock;
  assign CAMLine_39_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_39_io_wi = io_waddr[39]; // @[cam.scala 86:31]
  assign CAMLine_39_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_39_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_40_clock = clock;
  assign CAMLine_40_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_40_io_wi = io_waddr[40]; // @[cam.scala 86:31]
  assign CAMLine_40_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_40_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_41_clock = clock;
  assign CAMLine_41_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_41_io_wi = io_waddr[41]; // @[cam.scala 86:31]
  assign CAMLine_41_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_41_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_42_clock = clock;
  assign CAMLine_42_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_42_io_wi = io_waddr[42]; // @[cam.scala 86:31]
  assign CAMLine_42_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_42_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_43_clock = clock;
  assign CAMLine_43_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_43_io_wi = io_waddr[43]; // @[cam.scala 86:31]
  assign CAMLine_43_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_43_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_44_clock = clock;
  assign CAMLine_44_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_44_io_wi = io_waddr[44]; // @[cam.scala 86:31]
  assign CAMLine_44_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_44_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_45_clock = clock;
  assign CAMLine_45_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_45_io_wi = io_waddr[45]; // @[cam.scala 86:31]
  assign CAMLine_45_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_45_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_46_clock = clock;
  assign CAMLine_46_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_46_io_wi = io_waddr[46]; // @[cam.scala 86:31]
  assign CAMLine_46_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_46_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_47_clock = clock;
  assign CAMLine_47_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_47_io_wi = io_waddr[47]; // @[cam.scala 86:31]
  assign CAMLine_47_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_47_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_48_clock = clock;
  assign CAMLine_48_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_48_io_wi = io_waddr[48]; // @[cam.scala 86:31]
  assign CAMLine_48_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_48_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_49_clock = clock;
  assign CAMLine_49_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_49_io_wi = io_waddr[49]; // @[cam.scala 86:31]
  assign CAMLine_49_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_49_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_50_clock = clock;
  assign CAMLine_50_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_50_io_wi = io_waddr[50]; // @[cam.scala 86:31]
  assign CAMLine_50_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_50_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_51_clock = clock;
  assign CAMLine_51_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_51_io_wi = io_waddr[51]; // @[cam.scala 86:31]
  assign CAMLine_51_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_51_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_52_clock = clock;
  assign CAMLine_52_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_52_io_wi = io_waddr[52]; // @[cam.scala 86:31]
  assign CAMLine_52_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_52_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_53_clock = clock;
  assign CAMLine_53_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_53_io_wi = io_waddr[53]; // @[cam.scala 86:31]
  assign CAMLine_53_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_53_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_54_clock = clock;
  assign CAMLine_54_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_54_io_wi = io_waddr[54]; // @[cam.scala 86:31]
  assign CAMLine_54_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_54_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_55_clock = clock;
  assign CAMLine_55_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_55_io_wi = io_waddr[55]; // @[cam.scala 86:31]
  assign CAMLine_55_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_55_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_56_clock = clock;
  assign CAMLine_56_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_56_io_wi = io_waddr[56]; // @[cam.scala 86:31]
  assign CAMLine_56_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_56_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_57_clock = clock;
  assign CAMLine_57_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_57_io_wi = io_waddr[57]; // @[cam.scala 86:31]
  assign CAMLine_57_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_57_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_58_clock = clock;
  assign CAMLine_58_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_58_io_wi = io_waddr[58]; // @[cam.scala 86:31]
  assign CAMLine_58_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_58_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_59_clock = clock;
  assign CAMLine_59_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_59_io_wi = io_waddr[59]; // @[cam.scala 86:31]
  assign CAMLine_59_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_59_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_60_clock = clock;
  assign CAMLine_60_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_60_io_wi = io_waddr[60]; // @[cam.scala 86:31]
  assign CAMLine_60_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_60_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_61_clock = clock;
  assign CAMLine_61_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_61_io_wi = io_waddr[61]; // @[cam.scala 86:31]
  assign CAMLine_61_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_61_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_62_clock = clock;
  assign CAMLine_62_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_62_io_wi = io_waddr[62]; // @[cam.scala 86:31]
  assign CAMLine_62_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_62_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_63_clock = clock;
  assign CAMLine_63_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_63_io_wi = io_waddr[63]; // @[cam.scala 86:31]
  assign CAMLine_63_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_63_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_64_clock = clock;
  assign CAMLine_64_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_64_io_wi = io_waddr[64]; // @[cam.scala 86:31]
  assign CAMLine_64_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_64_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_65_clock = clock;
  assign CAMLine_65_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_65_io_wi = io_waddr[65]; // @[cam.scala 86:31]
  assign CAMLine_65_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_65_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_66_clock = clock;
  assign CAMLine_66_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_66_io_wi = io_waddr[66]; // @[cam.scala 86:31]
  assign CAMLine_66_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_66_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_67_clock = clock;
  assign CAMLine_67_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_67_io_wi = io_waddr[67]; // @[cam.scala 86:31]
  assign CAMLine_67_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_67_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_68_clock = clock;
  assign CAMLine_68_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_68_io_wi = io_waddr[68]; // @[cam.scala 86:31]
  assign CAMLine_68_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_68_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_69_clock = clock;
  assign CAMLine_69_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_69_io_wi = io_waddr[69]; // @[cam.scala 86:31]
  assign CAMLine_69_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_69_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_70_clock = clock;
  assign CAMLine_70_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_70_io_wi = io_waddr[70]; // @[cam.scala 86:31]
  assign CAMLine_70_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_70_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_71_clock = clock;
  assign CAMLine_71_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_71_io_wi = io_waddr[71]; // @[cam.scala 86:31]
  assign CAMLine_71_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_71_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_72_clock = clock;
  assign CAMLine_72_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_72_io_wi = io_waddr[72]; // @[cam.scala 86:31]
  assign CAMLine_72_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_72_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_73_clock = clock;
  assign CAMLine_73_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_73_io_wi = io_waddr[73]; // @[cam.scala 86:31]
  assign CAMLine_73_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_73_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_74_clock = clock;
  assign CAMLine_74_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_74_io_wi = io_waddr[74]; // @[cam.scala 86:31]
  assign CAMLine_74_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_74_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_75_clock = clock;
  assign CAMLine_75_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_75_io_wi = io_waddr[75]; // @[cam.scala 86:31]
  assign CAMLine_75_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_75_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_76_clock = clock;
  assign CAMLine_76_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_76_io_wi = io_waddr[76]; // @[cam.scala 86:31]
  assign CAMLine_76_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_76_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_77_clock = clock;
  assign CAMLine_77_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_77_io_wi = io_waddr[77]; // @[cam.scala 86:31]
  assign CAMLine_77_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_77_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_78_clock = clock;
  assign CAMLine_78_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_78_io_wi = io_waddr[78]; // @[cam.scala 86:31]
  assign CAMLine_78_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_78_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_79_clock = clock;
  assign CAMLine_79_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_79_io_wi = io_waddr[79]; // @[cam.scala 86:31]
  assign CAMLine_79_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_79_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_80_clock = clock;
  assign CAMLine_80_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_80_io_wi = io_waddr[80]; // @[cam.scala 86:31]
  assign CAMLine_80_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_80_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_81_clock = clock;
  assign CAMLine_81_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_81_io_wi = io_waddr[81]; // @[cam.scala 86:31]
  assign CAMLine_81_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_81_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_82_clock = clock;
  assign CAMLine_82_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_82_io_wi = io_waddr[82]; // @[cam.scala 86:31]
  assign CAMLine_82_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_82_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_83_clock = clock;
  assign CAMLine_83_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_83_io_wi = io_waddr[83]; // @[cam.scala 86:31]
  assign CAMLine_83_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_83_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_84_clock = clock;
  assign CAMLine_84_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_84_io_wi = io_waddr[84]; // @[cam.scala 86:31]
  assign CAMLine_84_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_84_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_85_clock = clock;
  assign CAMLine_85_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_85_io_wi = io_waddr[85]; // @[cam.scala 86:31]
  assign CAMLine_85_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_85_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_86_clock = clock;
  assign CAMLine_86_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_86_io_wi = io_waddr[86]; // @[cam.scala 86:31]
  assign CAMLine_86_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_86_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_87_clock = clock;
  assign CAMLine_87_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_87_io_wi = io_waddr[87]; // @[cam.scala 86:31]
  assign CAMLine_87_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_87_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_88_clock = clock;
  assign CAMLine_88_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_88_io_wi = io_waddr[88]; // @[cam.scala 86:31]
  assign CAMLine_88_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_88_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_89_clock = clock;
  assign CAMLine_89_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_89_io_wi = io_waddr[89]; // @[cam.scala 86:31]
  assign CAMLine_89_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_89_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_90_clock = clock;
  assign CAMLine_90_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_90_io_wi = io_waddr[90]; // @[cam.scala 86:31]
  assign CAMLine_90_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_90_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_91_clock = clock;
  assign CAMLine_91_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_91_io_wi = io_waddr[91]; // @[cam.scala 86:31]
  assign CAMLine_91_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_91_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_92_clock = clock;
  assign CAMLine_92_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_92_io_wi = io_waddr[92]; // @[cam.scala 86:31]
  assign CAMLine_92_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_92_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_93_clock = clock;
  assign CAMLine_93_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_93_io_wi = io_waddr[93]; // @[cam.scala 86:31]
  assign CAMLine_93_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_93_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_94_clock = clock;
  assign CAMLine_94_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_94_io_wi = io_waddr[94]; // @[cam.scala 86:31]
  assign CAMLine_94_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_94_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_95_clock = clock;
  assign CAMLine_95_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_95_io_wi = io_waddr[95]; // @[cam.scala 86:31]
  assign CAMLine_95_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_95_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_96_clock = clock;
  assign CAMLine_96_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_96_io_wi = io_waddr[96]; // @[cam.scala 86:31]
  assign CAMLine_96_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_96_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_97_clock = clock;
  assign CAMLine_97_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_97_io_wi = io_waddr[97]; // @[cam.scala 86:31]
  assign CAMLine_97_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_97_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_98_clock = clock;
  assign CAMLine_98_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_98_io_wi = io_waddr[98]; // @[cam.scala 86:31]
  assign CAMLine_98_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_98_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_99_clock = clock;
  assign CAMLine_99_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_99_io_wi = io_waddr[99]; // @[cam.scala 86:31]
  assign CAMLine_99_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_99_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_100_clock = clock;
  assign CAMLine_100_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_100_io_wi = io_waddr[100]; // @[cam.scala 86:31]
  assign CAMLine_100_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_100_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_101_clock = clock;
  assign CAMLine_101_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_101_io_wi = io_waddr[101]; // @[cam.scala 86:31]
  assign CAMLine_101_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_101_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_102_clock = clock;
  assign CAMLine_102_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_102_io_wi = io_waddr[102]; // @[cam.scala 86:31]
  assign CAMLine_102_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_102_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_103_clock = clock;
  assign CAMLine_103_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_103_io_wi = io_waddr[103]; // @[cam.scala 86:31]
  assign CAMLine_103_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_103_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_104_clock = clock;
  assign CAMLine_104_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_104_io_wi = io_waddr[104]; // @[cam.scala 86:31]
  assign CAMLine_104_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_104_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_105_clock = clock;
  assign CAMLine_105_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_105_io_wi = io_waddr[105]; // @[cam.scala 86:31]
  assign CAMLine_105_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_105_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_106_clock = clock;
  assign CAMLine_106_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_106_io_wi = io_waddr[106]; // @[cam.scala 86:31]
  assign CAMLine_106_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_106_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_107_clock = clock;
  assign CAMLine_107_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_107_io_wi = io_waddr[107]; // @[cam.scala 86:31]
  assign CAMLine_107_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_107_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_108_clock = clock;
  assign CAMLine_108_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_108_io_wi = io_waddr[108]; // @[cam.scala 86:31]
  assign CAMLine_108_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_108_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_109_clock = clock;
  assign CAMLine_109_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_109_io_wi = io_waddr[109]; // @[cam.scala 86:31]
  assign CAMLine_109_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_109_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_110_clock = clock;
  assign CAMLine_110_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_110_io_wi = io_waddr[110]; // @[cam.scala 86:31]
  assign CAMLine_110_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_110_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_111_clock = clock;
  assign CAMLine_111_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_111_io_wi = io_waddr[111]; // @[cam.scala 86:31]
  assign CAMLine_111_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_111_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_112_clock = clock;
  assign CAMLine_112_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_112_io_wi = io_waddr[112]; // @[cam.scala 86:31]
  assign CAMLine_112_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_112_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_113_clock = clock;
  assign CAMLine_113_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_113_io_wi = io_waddr[113]; // @[cam.scala 86:31]
  assign CAMLine_113_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_113_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_114_clock = clock;
  assign CAMLine_114_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_114_io_wi = io_waddr[114]; // @[cam.scala 86:31]
  assign CAMLine_114_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_114_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_115_clock = clock;
  assign CAMLine_115_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_115_io_wi = io_waddr[115]; // @[cam.scala 86:31]
  assign CAMLine_115_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_115_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_116_clock = clock;
  assign CAMLine_116_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_116_io_wi = io_waddr[116]; // @[cam.scala 86:31]
  assign CAMLine_116_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_116_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_117_clock = clock;
  assign CAMLine_117_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_117_io_wi = io_waddr[117]; // @[cam.scala 86:31]
  assign CAMLine_117_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_117_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_118_clock = clock;
  assign CAMLine_118_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_118_io_wi = io_waddr[118]; // @[cam.scala 86:31]
  assign CAMLine_118_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_118_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_119_clock = clock;
  assign CAMLine_119_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_119_io_wi = io_waddr[119]; // @[cam.scala 86:31]
  assign CAMLine_119_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_119_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_120_clock = clock;
  assign CAMLine_120_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_120_io_wi = io_waddr[120]; // @[cam.scala 86:31]
  assign CAMLine_120_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_120_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_121_clock = clock;
  assign CAMLine_121_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_121_io_wi = io_waddr[121]; // @[cam.scala 86:31]
  assign CAMLine_121_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_121_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_122_clock = clock;
  assign CAMLine_122_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_122_io_wi = io_waddr[122]; // @[cam.scala 86:31]
  assign CAMLine_122_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_122_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_123_clock = clock;
  assign CAMLine_123_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_123_io_wi = io_waddr[123]; // @[cam.scala 86:31]
  assign CAMLine_123_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_123_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_124_clock = clock;
  assign CAMLine_124_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_124_io_wi = io_waddr[124]; // @[cam.scala 86:31]
  assign CAMLine_124_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_124_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_125_clock = clock;
  assign CAMLine_125_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_125_io_wi = io_waddr[125]; // @[cam.scala 86:31]
  assign CAMLine_125_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_125_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_126_clock = clock;
  assign CAMLine_126_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_126_io_wi = io_waddr[126]; // @[cam.scala 86:31]
  assign CAMLine_126_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_126_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_127_clock = clock;
  assign CAMLine_127_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_127_io_wi = io_waddr[127]; // @[cam.scala 86:31]
  assign CAMLine_127_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_127_io_din = io_din; // @[cam.scala 88:21]
endmodule
