module FIFO(
  input          clock,
  input          reset,
  input          io_rst,
  input  [127:0] io_dataIn,
  input          io_push,
  input          io_pop,
  output [127:0] io_dataOut,
  output         io_full,
  output         io_empty
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [127:0] _RAND_27;
  reg [127:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [127:0] _RAND_33;
  reg [127:0] _RAND_34;
  reg [127:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [127:0] _RAND_38;
  reg [127:0] _RAND_39;
  reg [127:0] _RAND_40;
  reg [127:0] _RAND_41;
  reg [127:0] _RAND_42;
  reg [127:0] _RAND_43;
  reg [127:0] _RAND_44;
  reg [127:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [127:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [127:0] _RAND_50;
  reg [127:0] _RAND_51;
  reg [127:0] _RAND_52;
  reg [127:0] _RAND_53;
  reg [127:0] _RAND_54;
  reg [127:0] _RAND_55;
  reg [127:0] _RAND_56;
  reg [127:0] _RAND_57;
  reg [127:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [127:0] _RAND_61;
  reg [127:0] _RAND_62;
  reg [127:0] _RAND_63;
  reg [127:0] _RAND_64;
  reg [127:0] _RAND_65;
  reg [127:0] _RAND_66;
  reg [127:0] _RAND_67;
  reg [127:0] _RAND_68;
  reg [127:0] _RAND_69;
  reg [127:0] _RAND_70;
  reg [127:0] _RAND_71;
  reg [127:0] _RAND_72;
  reg [127:0] _RAND_73;
  reg [127:0] _RAND_74;
  reg [127:0] _RAND_75;
  reg [127:0] _RAND_76;
  reg [127:0] _RAND_77;
  reg [127:0] _RAND_78;
  reg [127:0] _RAND_79;
  reg [127:0] _RAND_80;
  reg [127:0] _RAND_81;
  reg [127:0] _RAND_82;
  reg [127:0] _RAND_83;
  reg [127:0] _RAND_84;
  reg [127:0] _RAND_85;
  reg [127:0] _RAND_86;
  reg [127:0] _RAND_87;
  reg [127:0] _RAND_88;
  reg [127:0] _RAND_89;
  reg [127:0] _RAND_90;
  reg [127:0] _RAND_91;
  reg [127:0] _RAND_92;
  reg [127:0] _RAND_93;
  reg [127:0] _RAND_94;
  reg [127:0] _RAND_95;
  reg [127:0] _RAND_96;
  reg [127:0] _RAND_97;
  reg [127:0] _RAND_98;
  reg [127:0] _RAND_99;
  reg [127:0] _RAND_100;
  reg [127:0] _RAND_101;
  reg [127:0] _RAND_102;
  reg [127:0] _RAND_103;
  reg [127:0] _RAND_104;
  reg [127:0] _RAND_105;
  reg [127:0] _RAND_106;
  reg [127:0] _RAND_107;
  reg [127:0] _RAND_108;
  reg [127:0] _RAND_109;
  reg [127:0] _RAND_110;
  reg [127:0] _RAND_111;
  reg [127:0] _RAND_112;
  reg [127:0] _RAND_113;
  reg [127:0] _RAND_114;
  reg [127:0] _RAND_115;
  reg [127:0] _RAND_116;
  reg [127:0] _RAND_117;
  reg [127:0] _RAND_118;
  reg [127:0] _RAND_119;
  reg [127:0] _RAND_120;
  reg [127:0] _RAND_121;
  reg [127:0] _RAND_122;
  reg [127:0] _RAND_123;
  reg [127:0] _RAND_124;
  reg [127:0] _RAND_125;
  reg [127:0] _RAND_126;
  reg [127:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] memRegs_0; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_1; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_2; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_3; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_4; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_5; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_6; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_7; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_8; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_9; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_10; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_11; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_12; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_13; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_14; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_15; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_16; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_17; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_18; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_19; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_20; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_21; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_22; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_23; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_24; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_25; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_26; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_27; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_28; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_29; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_30; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_31; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_32; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_33; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_34; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_35; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_36; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_37; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_38; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_39; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_40; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_41; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_42; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_43; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_44; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_45; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_46; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_47; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_48; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_49; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_50; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_51; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_52; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_53; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_54; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_55; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_56; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_57; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_58; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_59; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_60; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_61; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_62; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_63; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_64; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_65; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_66; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_67; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_68; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_69; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_70; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_71; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_72; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_73; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_74; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_75; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_76; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_77; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_78; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_79; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_80; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_81; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_82; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_83; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_84; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_85; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_86; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_87; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_88; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_89; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_90; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_91; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_92; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_93; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_94; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_95; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_96; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_97; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_98; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_99; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_100; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_101; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_102; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_103; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_104; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_105; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_106; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_107; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_108; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_109; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_110; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_111; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_112; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_113; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_114; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_115; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_116; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_117; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_118; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_119; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_120; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_121; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_122; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_123; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_124; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_125; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_126; // @[FIFO.scala 17:20]
  reg [127:0] memRegs_127; // @[FIFO.scala 17:20]
  reg [6:0] tailReg; // @[FIFO.scala 18:21]
  reg [6:0] headReg; // @[FIFO.scala 19:21]
  reg  emptyReg; // @[FIFO.scala 20:21]
  wire [6:0] _headReg_T_1 = headReg + 7'h1; // @[FIFO.scala 27:24]
  wire  _T_2 = ~emptyReg; // @[FIFO.scala 29:23]
  wire [6:0] _tailReg_T_1 = tailReg + 7'h1; // @[FIFO.scala 30:24]
  wire  _GEN_128 = _tailReg_T_1 == headReg | emptyReg; // @[FIFO.scala 31:39 32:16 20:21]
  wire  _GEN_130 = io_pop & ~emptyReg ? _GEN_128 : emptyReg; // @[FIFO.scala 20:21 29:34]
  wire  _GEN_260 = io_push & ~io_full ? 1'h0 : _GEN_130; // @[FIFO.scala 25:34 28:14]
  wire [127:0] _GEN_394 = 7'h1 == tailReg ? memRegs_1 : memRegs_0; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_395 = 7'h2 == tailReg ? memRegs_2 : _GEN_394; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_396 = 7'h3 == tailReg ? memRegs_3 : _GEN_395; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_397 = 7'h4 == tailReg ? memRegs_4 : _GEN_396; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_398 = 7'h5 == tailReg ? memRegs_5 : _GEN_397; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_399 = 7'h6 == tailReg ? memRegs_6 : _GEN_398; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_400 = 7'h7 == tailReg ? memRegs_7 : _GEN_399; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_401 = 7'h8 == tailReg ? memRegs_8 : _GEN_400; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_402 = 7'h9 == tailReg ? memRegs_9 : _GEN_401; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_403 = 7'ha == tailReg ? memRegs_10 : _GEN_402; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_404 = 7'hb == tailReg ? memRegs_11 : _GEN_403; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_405 = 7'hc == tailReg ? memRegs_12 : _GEN_404; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_406 = 7'hd == tailReg ? memRegs_13 : _GEN_405; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_407 = 7'he == tailReg ? memRegs_14 : _GEN_406; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_408 = 7'hf == tailReg ? memRegs_15 : _GEN_407; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_409 = 7'h10 == tailReg ? memRegs_16 : _GEN_408; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_410 = 7'h11 == tailReg ? memRegs_17 : _GEN_409; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_411 = 7'h12 == tailReg ? memRegs_18 : _GEN_410; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_412 = 7'h13 == tailReg ? memRegs_19 : _GEN_411; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_413 = 7'h14 == tailReg ? memRegs_20 : _GEN_412; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_414 = 7'h15 == tailReg ? memRegs_21 : _GEN_413; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_415 = 7'h16 == tailReg ? memRegs_22 : _GEN_414; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_416 = 7'h17 == tailReg ? memRegs_23 : _GEN_415; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_417 = 7'h18 == tailReg ? memRegs_24 : _GEN_416; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_418 = 7'h19 == tailReg ? memRegs_25 : _GEN_417; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_419 = 7'h1a == tailReg ? memRegs_26 : _GEN_418; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_420 = 7'h1b == tailReg ? memRegs_27 : _GEN_419; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_421 = 7'h1c == tailReg ? memRegs_28 : _GEN_420; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_422 = 7'h1d == tailReg ? memRegs_29 : _GEN_421; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_423 = 7'h1e == tailReg ? memRegs_30 : _GEN_422; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_424 = 7'h1f == tailReg ? memRegs_31 : _GEN_423; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_425 = 7'h20 == tailReg ? memRegs_32 : _GEN_424; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_426 = 7'h21 == tailReg ? memRegs_33 : _GEN_425; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_427 = 7'h22 == tailReg ? memRegs_34 : _GEN_426; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_428 = 7'h23 == tailReg ? memRegs_35 : _GEN_427; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_429 = 7'h24 == tailReg ? memRegs_36 : _GEN_428; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_430 = 7'h25 == tailReg ? memRegs_37 : _GEN_429; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_431 = 7'h26 == tailReg ? memRegs_38 : _GEN_430; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_432 = 7'h27 == tailReg ? memRegs_39 : _GEN_431; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_433 = 7'h28 == tailReg ? memRegs_40 : _GEN_432; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_434 = 7'h29 == tailReg ? memRegs_41 : _GEN_433; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_435 = 7'h2a == tailReg ? memRegs_42 : _GEN_434; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_436 = 7'h2b == tailReg ? memRegs_43 : _GEN_435; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_437 = 7'h2c == tailReg ? memRegs_44 : _GEN_436; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_438 = 7'h2d == tailReg ? memRegs_45 : _GEN_437; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_439 = 7'h2e == tailReg ? memRegs_46 : _GEN_438; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_440 = 7'h2f == tailReg ? memRegs_47 : _GEN_439; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_441 = 7'h30 == tailReg ? memRegs_48 : _GEN_440; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_442 = 7'h31 == tailReg ? memRegs_49 : _GEN_441; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_443 = 7'h32 == tailReg ? memRegs_50 : _GEN_442; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_444 = 7'h33 == tailReg ? memRegs_51 : _GEN_443; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_445 = 7'h34 == tailReg ? memRegs_52 : _GEN_444; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_446 = 7'h35 == tailReg ? memRegs_53 : _GEN_445; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_447 = 7'h36 == tailReg ? memRegs_54 : _GEN_446; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_448 = 7'h37 == tailReg ? memRegs_55 : _GEN_447; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_449 = 7'h38 == tailReg ? memRegs_56 : _GEN_448; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_450 = 7'h39 == tailReg ? memRegs_57 : _GEN_449; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_451 = 7'h3a == tailReg ? memRegs_58 : _GEN_450; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_452 = 7'h3b == tailReg ? memRegs_59 : _GEN_451; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_453 = 7'h3c == tailReg ? memRegs_60 : _GEN_452; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_454 = 7'h3d == tailReg ? memRegs_61 : _GEN_453; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_455 = 7'h3e == tailReg ? memRegs_62 : _GEN_454; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_456 = 7'h3f == tailReg ? memRegs_63 : _GEN_455; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_457 = 7'h40 == tailReg ? memRegs_64 : _GEN_456; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_458 = 7'h41 == tailReg ? memRegs_65 : _GEN_457; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_459 = 7'h42 == tailReg ? memRegs_66 : _GEN_458; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_460 = 7'h43 == tailReg ? memRegs_67 : _GEN_459; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_461 = 7'h44 == tailReg ? memRegs_68 : _GEN_460; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_462 = 7'h45 == tailReg ? memRegs_69 : _GEN_461; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_463 = 7'h46 == tailReg ? memRegs_70 : _GEN_462; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_464 = 7'h47 == tailReg ? memRegs_71 : _GEN_463; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_465 = 7'h48 == tailReg ? memRegs_72 : _GEN_464; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_466 = 7'h49 == tailReg ? memRegs_73 : _GEN_465; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_467 = 7'h4a == tailReg ? memRegs_74 : _GEN_466; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_468 = 7'h4b == tailReg ? memRegs_75 : _GEN_467; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_469 = 7'h4c == tailReg ? memRegs_76 : _GEN_468; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_470 = 7'h4d == tailReg ? memRegs_77 : _GEN_469; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_471 = 7'h4e == tailReg ? memRegs_78 : _GEN_470; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_472 = 7'h4f == tailReg ? memRegs_79 : _GEN_471; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_473 = 7'h50 == tailReg ? memRegs_80 : _GEN_472; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_474 = 7'h51 == tailReg ? memRegs_81 : _GEN_473; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_475 = 7'h52 == tailReg ? memRegs_82 : _GEN_474; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_476 = 7'h53 == tailReg ? memRegs_83 : _GEN_475; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_477 = 7'h54 == tailReg ? memRegs_84 : _GEN_476; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_478 = 7'h55 == tailReg ? memRegs_85 : _GEN_477; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_479 = 7'h56 == tailReg ? memRegs_86 : _GEN_478; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_480 = 7'h57 == tailReg ? memRegs_87 : _GEN_479; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_481 = 7'h58 == tailReg ? memRegs_88 : _GEN_480; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_482 = 7'h59 == tailReg ? memRegs_89 : _GEN_481; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_483 = 7'h5a == tailReg ? memRegs_90 : _GEN_482; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_484 = 7'h5b == tailReg ? memRegs_91 : _GEN_483; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_485 = 7'h5c == tailReg ? memRegs_92 : _GEN_484; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_486 = 7'h5d == tailReg ? memRegs_93 : _GEN_485; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_487 = 7'h5e == tailReg ? memRegs_94 : _GEN_486; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_488 = 7'h5f == tailReg ? memRegs_95 : _GEN_487; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_489 = 7'h60 == tailReg ? memRegs_96 : _GEN_488; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_490 = 7'h61 == tailReg ? memRegs_97 : _GEN_489; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_491 = 7'h62 == tailReg ? memRegs_98 : _GEN_490; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_492 = 7'h63 == tailReg ? memRegs_99 : _GEN_491; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_493 = 7'h64 == tailReg ? memRegs_100 : _GEN_492; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_494 = 7'h65 == tailReg ? memRegs_101 : _GEN_493; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_495 = 7'h66 == tailReg ? memRegs_102 : _GEN_494; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_496 = 7'h67 == tailReg ? memRegs_103 : _GEN_495; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_497 = 7'h68 == tailReg ? memRegs_104 : _GEN_496; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_498 = 7'h69 == tailReg ? memRegs_105 : _GEN_497; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_499 = 7'h6a == tailReg ? memRegs_106 : _GEN_498; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_500 = 7'h6b == tailReg ? memRegs_107 : _GEN_499; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_501 = 7'h6c == tailReg ? memRegs_108 : _GEN_500; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_502 = 7'h6d == tailReg ? memRegs_109 : _GEN_501; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_503 = 7'h6e == tailReg ? memRegs_110 : _GEN_502; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_504 = 7'h6f == tailReg ? memRegs_111 : _GEN_503; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_505 = 7'h70 == tailReg ? memRegs_112 : _GEN_504; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_506 = 7'h71 == tailReg ? memRegs_113 : _GEN_505; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_507 = 7'h72 == tailReg ? memRegs_114 : _GEN_506; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_508 = 7'h73 == tailReg ? memRegs_115 : _GEN_507; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_509 = 7'h74 == tailReg ? memRegs_116 : _GEN_508; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_510 = 7'h75 == tailReg ? memRegs_117 : _GEN_509; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_511 = 7'h76 == tailReg ? memRegs_118 : _GEN_510; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_512 = 7'h77 == tailReg ? memRegs_119 : _GEN_511; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_513 = 7'h78 == tailReg ? memRegs_120 : _GEN_512; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_514 = 7'h79 == tailReg ? memRegs_121 : _GEN_513; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_515 = 7'h7a == tailReg ? memRegs_122 : _GEN_514; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_516 = 7'h7b == tailReg ? memRegs_123 : _GEN_515; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_517 = 7'h7c == tailReg ? memRegs_124 : _GEN_516; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_518 = 7'h7d == tailReg ? memRegs_125 : _GEN_517; // @[FIFO.scala 36:{14,14}]
  wire [127:0] _GEN_519 = 7'h7e == tailReg ? memRegs_126 : _GEN_518; // @[FIFO.scala 36:{14,14}]
  assign io_dataOut = 7'h7f == tailReg ? memRegs_127 : _GEN_519; // @[FIFO.scala 36:{14,14}]
  assign io_full = tailReg == headReg & _T_2; // @[FIFO.scala 37:36]
  assign io_empty = emptyReg; // @[FIFO.scala 35:12]
  always @(posedge clock) begin
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h0 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_0 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h1 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_1 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h2 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_2 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h3 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_3 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h4 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_4 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h5 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_5 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h6 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_6 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h7 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_7 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h8 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_8 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h9 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_9 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'ha == headReg) begin // @[FIFO.scala 26:22]
          memRegs_10 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'hb == headReg) begin // @[FIFO.scala 26:22]
          memRegs_11 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'hc == headReg) begin // @[FIFO.scala 26:22]
          memRegs_12 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'hd == headReg) begin // @[FIFO.scala 26:22]
          memRegs_13 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'he == headReg) begin // @[FIFO.scala 26:22]
          memRegs_14 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'hf == headReg) begin // @[FIFO.scala 26:22]
          memRegs_15 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h10 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_16 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h11 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_17 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h12 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_18 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h13 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_19 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h14 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_20 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h15 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_21 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h16 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_22 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h17 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_23 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h18 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_24 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h19 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_25 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h1a == headReg) begin // @[FIFO.scala 26:22]
          memRegs_26 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h1b == headReg) begin // @[FIFO.scala 26:22]
          memRegs_27 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h1c == headReg) begin // @[FIFO.scala 26:22]
          memRegs_28 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h1d == headReg) begin // @[FIFO.scala 26:22]
          memRegs_29 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h1e == headReg) begin // @[FIFO.scala 26:22]
          memRegs_30 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h1f == headReg) begin // @[FIFO.scala 26:22]
          memRegs_31 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h20 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_32 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h21 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_33 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h22 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_34 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h23 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_35 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h24 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_36 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h25 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_37 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h26 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_38 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h27 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_39 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h28 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_40 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h29 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_41 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h2a == headReg) begin // @[FIFO.scala 26:22]
          memRegs_42 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h2b == headReg) begin // @[FIFO.scala 26:22]
          memRegs_43 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h2c == headReg) begin // @[FIFO.scala 26:22]
          memRegs_44 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h2d == headReg) begin // @[FIFO.scala 26:22]
          memRegs_45 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h2e == headReg) begin // @[FIFO.scala 26:22]
          memRegs_46 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h2f == headReg) begin // @[FIFO.scala 26:22]
          memRegs_47 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h30 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_48 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h31 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_49 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h32 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_50 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h33 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_51 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h34 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_52 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h35 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_53 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h36 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_54 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h37 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_55 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h38 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_56 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h39 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_57 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h3a == headReg) begin // @[FIFO.scala 26:22]
          memRegs_58 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h3b == headReg) begin // @[FIFO.scala 26:22]
          memRegs_59 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h3c == headReg) begin // @[FIFO.scala 26:22]
          memRegs_60 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h3d == headReg) begin // @[FIFO.scala 26:22]
          memRegs_61 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h3e == headReg) begin // @[FIFO.scala 26:22]
          memRegs_62 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h3f == headReg) begin // @[FIFO.scala 26:22]
          memRegs_63 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h40 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_64 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h41 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_65 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h42 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_66 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h43 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_67 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h44 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_68 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h45 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_69 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h46 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_70 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h47 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_71 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h48 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_72 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h49 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_73 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h4a == headReg) begin // @[FIFO.scala 26:22]
          memRegs_74 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h4b == headReg) begin // @[FIFO.scala 26:22]
          memRegs_75 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h4c == headReg) begin // @[FIFO.scala 26:22]
          memRegs_76 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h4d == headReg) begin // @[FIFO.scala 26:22]
          memRegs_77 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h4e == headReg) begin // @[FIFO.scala 26:22]
          memRegs_78 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h4f == headReg) begin // @[FIFO.scala 26:22]
          memRegs_79 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h50 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_80 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h51 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_81 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h52 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_82 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h53 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_83 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h54 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_84 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h55 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_85 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h56 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_86 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h57 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_87 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h58 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_88 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h59 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_89 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h5a == headReg) begin // @[FIFO.scala 26:22]
          memRegs_90 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h5b == headReg) begin // @[FIFO.scala 26:22]
          memRegs_91 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h5c == headReg) begin // @[FIFO.scala 26:22]
          memRegs_92 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h5d == headReg) begin // @[FIFO.scala 26:22]
          memRegs_93 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h5e == headReg) begin // @[FIFO.scala 26:22]
          memRegs_94 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h5f == headReg) begin // @[FIFO.scala 26:22]
          memRegs_95 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h60 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_96 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h61 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_97 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h62 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_98 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h63 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_99 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h64 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_100 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h65 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_101 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h66 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_102 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h67 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_103 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h68 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_104 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h69 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_105 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h6a == headReg) begin // @[FIFO.scala 26:22]
          memRegs_106 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h6b == headReg) begin // @[FIFO.scala 26:22]
          memRegs_107 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h6c == headReg) begin // @[FIFO.scala 26:22]
          memRegs_108 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h6d == headReg) begin // @[FIFO.scala 26:22]
          memRegs_109 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h6e == headReg) begin // @[FIFO.scala 26:22]
          memRegs_110 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h6f == headReg) begin // @[FIFO.scala 26:22]
          memRegs_111 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h70 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_112 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h71 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_113 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h72 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_114 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h73 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_115 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h74 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_116 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h75 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_117 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h76 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_118 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h77 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_119 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h78 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_120 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h79 == headReg) begin // @[FIFO.scala 26:22]
          memRegs_121 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h7a == headReg) begin // @[FIFO.scala 26:22]
          memRegs_122 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h7b == headReg) begin // @[FIFO.scala 26:22]
          memRegs_123 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h7c == headReg) begin // @[FIFO.scala 26:22]
          memRegs_124 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h7d == headReg) begin // @[FIFO.scala 26:22]
          memRegs_125 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h7e == headReg) begin // @[FIFO.scala 26:22]
          memRegs_126 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (!(io_rst)) begin // @[FIFO.scala 21:15]
      if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
        if (7'h7f == headReg) begin // @[FIFO.scala 26:22]
          memRegs_127 <= io_dataIn; // @[FIFO.scala 26:22]
        end
      end
    end
    if (io_rst) begin // @[FIFO.scala 21:15]
      tailReg <= 7'h0; // @[FIFO.scala 22:13]
    end else if (!(io_push & ~io_full)) begin // @[FIFO.scala 25:34]
      if (io_pop & ~emptyReg) begin // @[FIFO.scala 29:34]
        tailReg <= _tailReg_T_1; // @[FIFO.scala 30:13]
      end
    end
    if (io_rst) begin // @[FIFO.scala 21:15]
      headReg <= 7'h0; // @[FIFO.scala 23:13]
    end else if (io_push & ~io_full) begin // @[FIFO.scala 25:34]
      headReg <= _headReg_T_1; // @[FIFO.scala 27:13]
    end
    emptyReg <= io_rst | _GEN_260; // @[FIFO.scala 21:15 24:14]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  memRegs_0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  memRegs_1 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  memRegs_2 = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  memRegs_3 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  memRegs_4 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  memRegs_5 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  memRegs_6 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  memRegs_7 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  memRegs_8 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  memRegs_9 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  memRegs_10 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  memRegs_11 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  memRegs_12 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  memRegs_13 = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  memRegs_14 = _RAND_14[127:0];
  _RAND_15 = {4{`RANDOM}};
  memRegs_15 = _RAND_15[127:0];
  _RAND_16 = {4{`RANDOM}};
  memRegs_16 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  memRegs_17 = _RAND_17[127:0];
  _RAND_18 = {4{`RANDOM}};
  memRegs_18 = _RAND_18[127:0];
  _RAND_19 = {4{`RANDOM}};
  memRegs_19 = _RAND_19[127:0];
  _RAND_20 = {4{`RANDOM}};
  memRegs_20 = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  memRegs_21 = _RAND_21[127:0];
  _RAND_22 = {4{`RANDOM}};
  memRegs_22 = _RAND_22[127:0];
  _RAND_23 = {4{`RANDOM}};
  memRegs_23 = _RAND_23[127:0];
  _RAND_24 = {4{`RANDOM}};
  memRegs_24 = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  memRegs_25 = _RAND_25[127:0];
  _RAND_26 = {4{`RANDOM}};
  memRegs_26 = _RAND_26[127:0];
  _RAND_27 = {4{`RANDOM}};
  memRegs_27 = _RAND_27[127:0];
  _RAND_28 = {4{`RANDOM}};
  memRegs_28 = _RAND_28[127:0];
  _RAND_29 = {4{`RANDOM}};
  memRegs_29 = _RAND_29[127:0];
  _RAND_30 = {4{`RANDOM}};
  memRegs_30 = _RAND_30[127:0];
  _RAND_31 = {4{`RANDOM}};
  memRegs_31 = _RAND_31[127:0];
  _RAND_32 = {4{`RANDOM}};
  memRegs_32 = _RAND_32[127:0];
  _RAND_33 = {4{`RANDOM}};
  memRegs_33 = _RAND_33[127:0];
  _RAND_34 = {4{`RANDOM}};
  memRegs_34 = _RAND_34[127:0];
  _RAND_35 = {4{`RANDOM}};
  memRegs_35 = _RAND_35[127:0];
  _RAND_36 = {4{`RANDOM}};
  memRegs_36 = _RAND_36[127:0];
  _RAND_37 = {4{`RANDOM}};
  memRegs_37 = _RAND_37[127:0];
  _RAND_38 = {4{`RANDOM}};
  memRegs_38 = _RAND_38[127:0];
  _RAND_39 = {4{`RANDOM}};
  memRegs_39 = _RAND_39[127:0];
  _RAND_40 = {4{`RANDOM}};
  memRegs_40 = _RAND_40[127:0];
  _RAND_41 = {4{`RANDOM}};
  memRegs_41 = _RAND_41[127:0];
  _RAND_42 = {4{`RANDOM}};
  memRegs_42 = _RAND_42[127:0];
  _RAND_43 = {4{`RANDOM}};
  memRegs_43 = _RAND_43[127:0];
  _RAND_44 = {4{`RANDOM}};
  memRegs_44 = _RAND_44[127:0];
  _RAND_45 = {4{`RANDOM}};
  memRegs_45 = _RAND_45[127:0];
  _RAND_46 = {4{`RANDOM}};
  memRegs_46 = _RAND_46[127:0];
  _RAND_47 = {4{`RANDOM}};
  memRegs_47 = _RAND_47[127:0];
  _RAND_48 = {4{`RANDOM}};
  memRegs_48 = _RAND_48[127:0];
  _RAND_49 = {4{`RANDOM}};
  memRegs_49 = _RAND_49[127:0];
  _RAND_50 = {4{`RANDOM}};
  memRegs_50 = _RAND_50[127:0];
  _RAND_51 = {4{`RANDOM}};
  memRegs_51 = _RAND_51[127:0];
  _RAND_52 = {4{`RANDOM}};
  memRegs_52 = _RAND_52[127:0];
  _RAND_53 = {4{`RANDOM}};
  memRegs_53 = _RAND_53[127:0];
  _RAND_54 = {4{`RANDOM}};
  memRegs_54 = _RAND_54[127:0];
  _RAND_55 = {4{`RANDOM}};
  memRegs_55 = _RAND_55[127:0];
  _RAND_56 = {4{`RANDOM}};
  memRegs_56 = _RAND_56[127:0];
  _RAND_57 = {4{`RANDOM}};
  memRegs_57 = _RAND_57[127:0];
  _RAND_58 = {4{`RANDOM}};
  memRegs_58 = _RAND_58[127:0];
  _RAND_59 = {4{`RANDOM}};
  memRegs_59 = _RAND_59[127:0];
  _RAND_60 = {4{`RANDOM}};
  memRegs_60 = _RAND_60[127:0];
  _RAND_61 = {4{`RANDOM}};
  memRegs_61 = _RAND_61[127:0];
  _RAND_62 = {4{`RANDOM}};
  memRegs_62 = _RAND_62[127:0];
  _RAND_63 = {4{`RANDOM}};
  memRegs_63 = _RAND_63[127:0];
  _RAND_64 = {4{`RANDOM}};
  memRegs_64 = _RAND_64[127:0];
  _RAND_65 = {4{`RANDOM}};
  memRegs_65 = _RAND_65[127:0];
  _RAND_66 = {4{`RANDOM}};
  memRegs_66 = _RAND_66[127:0];
  _RAND_67 = {4{`RANDOM}};
  memRegs_67 = _RAND_67[127:0];
  _RAND_68 = {4{`RANDOM}};
  memRegs_68 = _RAND_68[127:0];
  _RAND_69 = {4{`RANDOM}};
  memRegs_69 = _RAND_69[127:0];
  _RAND_70 = {4{`RANDOM}};
  memRegs_70 = _RAND_70[127:0];
  _RAND_71 = {4{`RANDOM}};
  memRegs_71 = _RAND_71[127:0];
  _RAND_72 = {4{`RANDOM}};
  memRegs_72 = _RAND_72[127:0];
  _RAND_73 = {4{`RANDOM}};
  memRegs_73 = _RAND_73[127:0];
  _RAND_74 = {4{`RANDOM}};
  memRegs_74 = _RAND_74[127:0];
  _RAND_75 = {4{`RANDOM}};
  memRegs_75 = _RAND_75[127:0];
  _RAND_76 = {4{`RANDOM}};
  memRegs_76 = _RAND_76[127:0];
  _RAND_77 = {4{`RANDOM}};
  memRegs_77 = _RAND_77[127:0];
  _RAND_78 = {4{`RANDOM}};
  memRegs_78 = _RAND_78[127:0];
  _RAND_79 = {4{`RANDOM}};
  memRegs_79 = _RAND_79[127:0];
  _RAND_80 = {4{`RANDOM}};
  memRegs_80 = _RAND_80[127:0];
  _RAND_81 = {4{`RANDOM}};
  memRegs_81 = _RAND_81[127:0];
  _RAND_82 = {4{`RANDOM}};
  memRegs_82 = _RAND_82[127:0];
  _RAND_83 = {4{`RANDOM}};
  memRegs_83 = _RAND_83[127:0];
  _RAND_84 = {4{`RANDOM}};
  memRegs_84 = _RAND_84[127:0];
  _RAND_85 = {4{`RANDOM}};
  memRegs_85 = _RAND_85[127:0];
  _RAND_86 = {4{`RANDOM}};
  memRegs_86 = _RAND_86[127:0];
  _RAND_87 = {4{`RANDOM}};
  memRegs_87 = _RAND_87[127:0];
  _RAND_88 = {4{`RANDOM}};
  memRegs_88 = _RAND_88[127:0];
  _RAND_89 = {4{`RANDOM}};
  memRegs_89 = _RAND_89[127:0];
  _RAND_90 = {4{`RANDOM}};
  memRegs_90 = _RAND_90[127:0];
  _RAND_91 = {4{`RANDOM}};
  memRegs_91 = _RAND_91[127:0];
  _RAND_92 = {4{`RANDOM}};
  memRegs_92 = _RAND_92[127:0];
  _RAND_93 = {4{`RANDOM}};
  memRegs_93 = _RAND_93[127:0];
  _RAND_94 = {4{`RANDOM}};
  memRegs_94 = _RAND_94[127:0];
  _RAND_95 = {4{`RANDOM}};
  memRegs_95 = _RAND_95[127:0];
  _RAND_96 = {4{`RANDOM}};
  memRegs_96 = _RAND_96[127:0];
  _RAND_97 = {4{`RANDOM}};
  memRegs_97 = _RAND_97[127:0];
  _RAND_98 = {4{`RANDOM}};
  memRegs_98 = _RAND_98[127:0];
  _RAND_99 = {4{`RANDOM}};
  memRegs_99 = _RAND_99[127:0];
  _RAND_100 = {4{`RANDOM}};
  memRegs_100 = _RAND_100[127:0];
  _RAND_101 = {4{`RANDOM}};
  memRegs_101 = _RAND_101[127:0];
  _RAND_102 = {4{`RANDOM}};
  memRegs_102 = _RAND_102[127:0];
  _RAND_103 = {4{`RANDOM}};
  memRegs_103 = _RAND_103[127:0];
  _RAND_104 = {4{`RANDOM}};
  memRegs_104 = _RAND_104[127:0];
  _RAND_105 = {4{`RANDOM}};
  memRegs_105 = _RAND_105[127:0];
  _RAND_106 = {4{`RANDOM}};
  memRegs_106 = _RAND_106[127:0];
  _RAND_107 = {4{`RANDOM}};
  memRegs_107 = _RAND_107[127:0];
  _RAND_108 = {4{`RANDOM}};
  memRegs_108 = _RAND_108[127:0];
  _RAND_109 = {4{`RANDOM}};
  memRegs_109 = _RAND_109[127:0];
  _RAND_110 = {4{`RANDOM}};
  memRegs_110 = _RAND_110[127:0];
  _RAND_111 = {4{`RANDOM}};
  memRegs_111 = _RAND_111[127:0];
  _RAND_112 = {4{`RANDOM}};
  memRegs_112 = _RAND_112[127:0];
  _RAND_113 = {4{`RANDOM}};
  memRegs_113 = _RAND_113[127:0];
  _RAND_114 = {4{`RANDOM}};
  memRegs_114 = _RAND_114[127:0];
  _RAND_115 = {4{`RANDOM}};
  memRegs_115 = _RAND_115[127:0];
  _RAND_116 = {4{`RANDOM}};
  memRegs_116 = _RAND_116[127:0];
  _RAND_117 = {4{`RANDOM}};
  memRegs_117 = _RAND_117[127:0];
  _RAND_118 = {4{`RANDOM}};
  memRegs_118 = _RAND_118[127:0];
  _RAND_119 = {4{`RANDOM}};
  memRegs_119 = _RAND_119[127:0];
  _RAND_120 = {4{`RANDOM}};
  memRegs_120 = _RAND_120[127:0];
  _RAND_121 = {4{`RANDOM}};
  memRegs_121 = _RAND_121[127:0];
  _RAND_122 = {4{`RANDOM}};
  memRegs_122 = _RAND_122[127:0];
  _RAND_123 = {4{`RANDOM}};
  memRegs_123 = _RAND_123[127:0];
  _RAND_124 = {4{`RANDOM}};
  memRegs_124 = _RAND_124[127:0];
  _RAND_125 = {4{`RANDOM}};
  memRegs_125 = _RAND_125[127:0];
  _RAND_126 = {4{`RANDOM}};
  memRegs_126 = _RAND_126[127:0];
  _RAND_127 = {4{`RANDOM}};
  memRegs_127 = _RAND_127[127:0];
  _RAND_128 = {1{`RANDOM}};
  tailReg = _RAND_128[6:0];
  _RAND_129 = {1{`RANDOM}};
  headReg = _RAND_129[6:0];
  _RAND_130 = {1{`RANDOM}};
  emptyReg = _RAND_130[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
