module Risc(
  input         clock,
  input         reset,
  input         io_isWr,
  input  [7:0]  io_wrAddr,
  input  [31:0] io_wrData,
  input         io_boot,
  output        io_valid,
  output [31:0] io_out
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] file [0:255]; // @[Risc.scala 16:17]
  wire  file_ra_MPORT_en; // @[Risc.scala 16:17]
  wire [7:0] file_ra_MPORT_addr; // @[Risc.scala 16:17]
  wire [31:0] file_ra_MPORT_data; // @[Risc.scala 16:17]
  wire  file_rb_MPORT_en; // @[Risc.scala 16:17]
  wire [7:0] file_rb_MPORT_addr; // @[Risc.scala 16:17]
  wire [31:0] file_rb_MPORT_data; // @[Risc.scala 16:17]
  wire [31:0] file_MPORT_data; // @[Risc.scala 16:17]
  wire [7:0] file_MPORT_addr; // @[Risc.scala 16:17]
  wire  file_MPORT_mask; // @[Risc.scala 16:17]
  wire  file_MPORT_en; // @[Risc.scala 16:17]
  reg [31:0] code_0; // @[Risc.scala 19:21]
  reg [31:0] code_1; // @[Risc.scala 19:21]
  reg [31:0] code_2; // @[Risc.scala 19:21]
  reg [31:0] code_3; // @[Risc.scala 19:21]
  reg [31:0] code_4; // @[Risc.scala 19:21]
  reg [31:0] code_5; // @[Risc.scala 19:21]
  reg [31:0] code_6; // @[Risc.scala 19:21]
  reg [31:0] code_7; // @[Risc.scala 19:21]
  reg [31:0] code_8; // @[Risc.scala 19:21]
  reg [31:0] code_9; // @[Risc.scala 19:21]
  reg [31:0] code_10; // @[Risc.scala 19:21]
  reg [31:0] code_11; // @[Risc.scala 19:21]
  reg [31:0] code_12; // @[Risc.scala 19:21]
  reg [31:0] code_13; // @[Risc.scala 19:21]
  reg [31:0] code_14; // @[Risc.scala 19:21]
  reg [31:0] code_15; // @[Risc.scala 19:21]
  reg [31:0] code_16; // @[Risc.scala 19:21]
  reg [31:0] code_17; // @[Risc.scala 19:21]
  reg [31:0] code_18; // @[Risc.scala 19:21]
  reg [31:0] code_19; // @[Risc.scala 19:21]
  reg [31:0] code_20; // @[Risc.scala 19:21]
  reg [31:0] code_21; // @[Risc.scala 19:21]
  reg [31:0] code_22; // @[Risc.scala 19:21]
  reg [31:0] code_23; // @[Risc.scala 19:21]
  reg [31:0] code_24; // @[Risc.scala 19:21]
  reg [31:0] code_25; // @[Risc.scala 19:21]
  reg [31:0] code_26; // @[Risc.scala 19:21]
  reg [31:0] code_27; // @[Risc.scala 19:21]
  reg [31:0] code_28; // @[Risc.scala 19:21]
  reg [31:0] code_29; // @[Risc.scala 19:21]
  reg [31:0] code_30; // @[Risc.scala 19:21]
  reg [31:0] code_31; // @[Risc.scala 19:21]
  reg [31:0] code_32; // @[Risc.scala 19:21]
  reg [31:0] code_33; // @[Risc.scala 19:21]
  reg [31:0] code_34; // @[Risc.scala 19:21]
  reg [31:0] code_35; // @[Risc.scala 19:21]
  reg [31:0] code_36; // @[Risc.scala 19:21]
  reg [31:0] code_37; // @[Risc.scala 19:21]
  reg [31:0] code_38; // @[Risc.scala 19:21]
  reg [31:0] code_39; // @[Risc.scala 19:21]
  reg [31:0] code_40; // @[Risc.scala 19:21]
  reg [31:0] code_41; // @[Risc.scala 19:21]
  reg [31:0] code_42; // @[Risc.scala 19:21]
  reg [31:0] code_43; // @[Risc.scala 19:21]
  reg [31:0] code_44; // @[Risc.scala 19:21]
  reg [31:0] code_45; // @[Risc.scala 19:21]
  reg [31:0] code_46; // @[Risc.scala 19:21]
  reg [31:0] code_47; // @[Risc.scala 19:21]
  reg [31:0] code_48; // @[Risc.scala 19:21]
  reg [31:0] code_49; // @[Risc.scala 19:21]
  reg [31:0] code_50; // @[Risc.scala 19:21]
  reg [31:0] code_51; // @[Risc.scala 19:21]
  reg [31:0] code_52; // @[Risc.scala 19:21]
  reg [31:0] code_53; // @[Risc.scala 19:21]
  reg [31:0] code_54; // @[Risc.scala 19:21]
  reg [31:0] code_55; // @[Risc.scala 19:21]
  reg [31:0] code_56; // @[Risc.scala 19:21]
  reg [31:0] code_57; // @[Risc.scala 19:21]
  reg [31:0] code_58; // @[Risc.scala 19:21]
  reg [31:0] code_59; // @[Risc.scala 19:21]
  reg [31:0] code_60; // @[Risc.scala 19:21]
  reg [31:0] code_61; // @[Risc.scala 19:21]
  reg [31:0] code_62; // @[Risc.scala 19:21]
  reg [31:0] code_63; // @[Risc.scala 19:21]
  reg [31:0] code_64; // @[Risc.scala 19:21]
  reg [31:0] code_65; // @[Risc.scala 19:21]
  reg [31:0] code_66; // @[Risc.scala 19:21]
  reg [31:0] code_67; // @[Risc.scala 19:21]
  reg [31:0] code_68; // @[Risc.scala 19:21]
  reg [31:0] code_69; // @[Risc.scala 19:21]
  reg [31:0] code_70; // @[Risc.scala 19:21]
  reg [31:0] code_71; // @[Risc.scala 19:21]
  reg [31:0] code_72; // @[Risc.scala 19:21]
  reg [31:0] code_73; // @[Risc.scala 19:21]
  reg [31:0] code_74; // @[Risc.scala 19:21]
  reg [31:0] code_75; // @[Risc.scala 19:21]
  reg [31:0] code_76; // @[Risc.scala 19:21]
  reg [31:0] code_77; // @[Risc.scala 19:21]
  reg [31:0] code_78; // @[Risc.scala 19:21]
  reg [31:0] code_79; // @[Risc.scala 19:21]
  reg [31:0] code_80; // @[Risc.scala 19:21]
  reg [31:0] code_81; // @[Risc.scala 19:21]
  reg [31:0] code_82; // @[Risc.scala 19:21]
  reg [31:0] code_83; // @[Risc.scala 19:21]
  reg [31:0] code_84; // @[Risc.scala 19:21]
  reg [31:0] code_85; // @[Risc.scala 19:21]
  reg [31:0] code_86; // @[Risc.scala 19:21]
  reg [31:0] code_87; // @[Risc.scala 19:21]
  reg [31:0] code_88; // @[Risc.scala 19:21]
  reg [31:0] code_89; // @[Risc.scala 19:21]
  reg [31:0] code_90; // @[Risc.scala 19:21]
  reg [31:0] code_91; // @[Risc.scala 19:21]
  reg [31:0] code_92; // @[Risc.scala 19:21]
  reg [31:0] code_93; // @[Risc.scala 19:21]
  reg [31:0] code_94; // @[Risc.scala 19:21]
  reg [31:0] code_95; // @[Risc.scala 19:21]
  reg [31:0] code_96; // @[Risc.scala 19:21]
  reg [31:0] code_97; // @[Risc.scala 19:21]
  reg [31:0] code_98; // @[Risc.scala 19:21]
  reg [31:0] code_99; // @[Risc.scala 19:21]
  reg [31:0] code_100; // @[Risc.scala 19:21]
  reg [31:0] code_101; // @[Risc.scala 19:21]
  reg [31:0] code_102; // @[Risc.scala 19:21]
  reg [31:0] code_103; // @[Risc.scala 19:21]
  reg [31:0] code_104; // @[Risc.scala 19:21]
  reg [31:0] code_105; // @[Risc.scala 19:21]
  reg [31:0] code_106; // @[Risc.scala 19:21]
  reg [31:0] code_107; // @[Risc.scala 19:21]
  reg [31:0] code_108; // @[Risc.scala 19:21]
  reg [31:0] code_109; // @[Risc.scala 19:21]
  reg [31:0] code_110; // @[Risc.scala 19:21]
  reg [31:0] code_111; // @[Risc.scala 19:21]
  reg [31:0] code_112; // @[Risc.scala 19:21]
  reg [31:0] code_113; // @[Risc.scala 19:21]
  reg [31:0] code_114; // @[Risc.scala 19:21]
  reg [31:0] code_115; // @[Risc.scala 19:21]
  reg [31:0] code_116; // @[Risc.scala 19:21]
  reg [31:0] code_117; // @[Risc.scala 19:21]
  reg [31:0] code_118; // @[Risc.scala 19:21]
  reg [31:0] code_119; // @[Risc.scala 19:21]
  reg [31:0] code_120; // @[Risc.scala 19:21]
  reg [31:0] code_121; // @[Risc.scala 19:21]
  reg [31:0] code_122; // @[Risc.scala 19:21]
  reg [31:0] code_123; // @[Risc.scala 19:21]
  reg [31:0] code_124; // @[Risc.scala 19:21]
  reg [31:0] code_125; // @[Risc.scala 19:21]
  reg [31:0] code_126; // @[Risc.scala 19:21]
  reg [31:0] code_127; // @[Risc.scala 19:21]
  reg [31:0] code_128; // @[Risc.scala 19:21]
  reg [31:0] code_129; // @[Risc.scala 19:21]
  reg [31:0] code_130; // @[Risc.scala 19:21]
  reg [31:0] code_131; // @[Risc.scala 19:21]
  reg [31:0] code_132; // @[Risc.scala 19:21]
  reg [31:0] code_133; // @[Risc.scala 19:21]
  reg [31:0] code_134; // @[Risc.scala 19:21]
  reg [31:0] code_135; // @[Risc.scala 19:21]
  reg [31:0] code_136; // @[Risc.scala 19:21]
  reg [31:0] code_137; // @[Risc.scala 19:21]
  reg [31:0] code_138; // @[Risc.scala 19:21]
  reg [31:0] code_139; // @[Risc.scala 19:21]
  reg [31:0] code_140; // @[Risc.scala 19:21]
  reg [31:0] code_141; // @[Risc.scala 19:21]
  reg [31:0] code_142; // @[Risc.scala 19:21]
  reg [31:0] code_143; // @[Risc.scala 19:21]
  reg [31:0] code_144; // @[Risc.scala 19:21]
  reg [31:0] code_145; // @[Risc.scala 19:21]
  reg [31:0] code_146; // @[Risc.scala 19:21]
  reg [31:0] code_147; // @[Risc.scala 19:21]
  reg [31:0] code_148; // @[Risc.scala 19:21]
  reg [31:0] code_149; // @[Risc.scala 19:21]
  reg [31:0] code_150; // @[Risc.scala 19:21]
  reg [31:0] code_151; // @[Risc.scala 19:21]
  reg [31:0] code_152; // @[Risc.scala 19:21]
  reg [31:0] code_153; // @[Risc.scala 19:21]
  reg [31:0] code_154; // @[Risc.scala 19:21]
  reg [31:0] code_155; // @[Risc.scala 19:21]
  reg [31:0] code_156; // @[Risc.scala 19:21]
  reg [31:0] code_157; // @[Risc.scala 19:21]
  reg [31:0] code_158; // @[Risc.scala 19:21]
  reg [31:0] code_159; // @[Risc.scala 19:21]
  reg [31:0] code_160; // @[Risc.scala 19:21]
  reg [31:0] code_161; // @[Risc.scala 19:21]
  reg [31:0] code_162; // @[Risc.scala 19:21]
  reg [31:0] code_163; // @[Risc.scala 19:21]
  reg [31:0] code_164; // @[Risc.scala 19:21]
  reg [31:0] code_165; // @[Risc.scala 19:21]
  reg [31:0] code_166; // @[Risc.scala 19:21]
  reg [31:0] code_167; // @[Risc.scala 19:21]
  reg [31:0] code_168; // @[Risc.scala 19:21]
  reg [31:0] code_169; // @[Risc.scala 19:21]
  reg [31:0] code_170; // @[Risc.scala 19:21]
  reg [31:0] code_171; // @[Risc.scala 19:21]
  reg [31:0] code_172; // @[Risc.scala 19:21]
  reg [31:0] code_173; // @[Risc.scala 19:21]
  reg [31:0] code_174; // @[Risc.scala 19:21]
  reg [31:0] code_175; // @[Risc.scala 19:21]
  reg [31:0] code_176; // @[Risc.scala 19:21]
  reg [31:0] code_177; // @[Risc.scala 19:21]
  reg [31:0] code_178; // @[Risc.scala 19:21]
  reg [31:0] code_179; // @[Risc.scala 19:21]
  reg [31:0] code_180; // @[Risc.scala 19:21]
  reg [31:0] code_181; // @[Risc.scala 19:21]
  reg [31:0] code_182; // @[Risc.scala 19:21]
  reg [31:0] code_183; // @[Risc.scala 19:21]
  reg [31:0] code_184; // @[Risc.scala 19:21]
  reg [31:0] code_185; // @[Risc.scala 19:21]
  reg [31:0] code_186; // @[Risc.scala 19:21]
  reg [31:0] code_187; // @[Risc.scala 19:21]
  reg [31:0] code_188; // @[Risc.scala 19:21]
  reg [31:0] code_189; // @[Risc.scala 19:21]
  reg [31:0] code_190; // @[Risc.scala 19:21]
  reg [31:0] code_191; // @[Risc.scala 19:21]
  reg [31:0] code_192; // @[Risc.scala 19:21]
  reg [31:0] code_193; // @[Risc.scala 19:21]
  reg [31:0] code_194; // @[Risc.scala 19:21]
  reg [31:0] code_195; // @[Risc.scala 19:21]
  reg [31:0] code_196; // @[Risc.scala 19:21]
  reg [31:0] code_197; // @[Risc.scala 19:21]
  reg [31:0] code_198; // @[Risc.scala 19:21]
  reg [31:0] code_199; // @[Risc.scala 19:21]
  reg [31:0] code_200; // @[Risc.scala 19:21]
  reg [31:0] code_201; // @[Risc.scala 19:21]
  reg [31:0] code_202; // @[Risc.scala 19:21]
  reg [31:0] code_203; // @[Risc.scala 19:21]
  reg [31:0] code_204; // @[Risc.scala 19:21]
  reg [31:0] code_205; // @[Risc.scala 19:21]
  reg [31:0] code_206; // @[Risc.scala 19:21]
  reg [31:0] code_207; // @[Risc.scala 19:21]
  reg [31:0] code_208; // @[Risc.scala 19:21]
  reg [31:0] code_209; // @[Risc.scala 19:21]
  reg [31:0] code_210; // @[Risc.scala 19:21]
  reg [31:0] code_211; // @[Risc.scala 19:21]
  reg [31:0] code_212; // @[Risc.scala 19:21]
  reg [31:0] code_213; // @[Risc.scala 19:21]
  reg [31:0] code_214; // @[Risc.scala 19:21]
  reg [31:0] code_215; // @[Risc.scala 19:21]
  reg [31:0] code_216; // @[Risc.scala 19:21]
  reg [31:0] code_217; // @[Risc.scala 19:21]
  reg [31:0] code_218; // @[Risc.scala 19:21]
  reg [31:0] code_219; // @[Risc.scala 19:21]
  reg [31:0] code_220; // @[Risc.scala 19:21]
  reg [31:0] code_221; // @[Risc.scala 19:21]
  reg [31:0] code_222; // @[Risc.scala 19:21]
  reg [31:0] code_223; // @[Risc.scala 19:21]
  reg [31:0] code_224; // @[Risc.scala 19:21]
  reg [31:0] code_225; // @[Risc.scala 19:21]
  reg [31:0] code_226; // @[Risc.scala 19:21]
  reg [31:0] code_227; // @[Risc.scala 19:21]
  reg [31:0] code_228; // @[Risc.scala 19:21]
  reg [31:0] code_229; // @[Risc.scala 19:21]
  reg [31:0] code_230; // @[Risc.scala 19:21]
  reg [31:0] code_231; // @[Risc.scala 19:21]
  reg [31:0] code_232; // @[Risc.scala 19:21]
  reg [31:0] code_233; // @[Risc.scala 19:21]
  reg [31:0] code_234; // @[Risc.scala 19:21]
  reg [31:0] code_235; // @[Risc.scala 19:21]
  reg [31:0] code_236; // @[Risc.scala 19:21]
  reg [31:0] code_237; // @[Risc.scala 19:21]
  reg [31:0] code_238; // @[Risc.scala 19:21]
  reg [31:0] code_239; // @[Risc.scala 19:21]
  reg [31:0] code_240; // @[Risc.scala 19:21]
  reg [31:0] code_241; // @[Risc.scala 19:21]
  reg [31:0] code_242; // @[Risc.scala 19:21]
  reg [31:0] code_243; // @[Risc.scala 19:21]
  reg [31:0] code_244; // @[Risc.scala 19:21]
  reg [31:0] code_245; // @[Risc.scala 19:21]
  reg [31:0] code_246; // @[Risc.scala 19:21]
  reg [31:0] code_247; // @[Risc.scala 19:21]
  reg [31:0] code_248; // @[Risc.scala 19:21]
  reg [31:0] code_249; // @[Risc.scala 19:21]
  reg [31:0] code_250; // @[Risc.scala 19:21]
  reg [31:0] code_251; // @[Risc.scala 19:21]
  reg [31:0] code_252; // @[Risc.scala 19:21]
  reg [31:0] code_253; // @[Risc.scala 19:21]
  reg [31:0] code_254; // @[Risc.scala 19:21]
  reg [31:0] code_255; // @[Risc.scala 19:21]
  reg [7:0] pc; // @[Risc.scala 21:21]
  wire [31:0] _GEN_1 = 8'h1 == pc ? code_1 : code_0; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_2 = 8'h2 == pc ? code_2 : _GEN_1; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_3 = 8'h3 == pc ? code_3 : _GEN_2; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_4 = 8'h4 == pc ? code_4 : _GEN_3; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_5 = 8'h5 == pc ? code_5 : _GEN_4; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_6 = 8'h6 == pc ? code_6 : _GEN_5; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_7 = 8'h7 == pc ? code_7 : _GEN_6; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_8 = 8'h8 == pc ? code_8 : _GEN_7; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_9 = 8'h9 == pc ? code_9 : _GEN_8; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_10 = 8'ha == pc ? code_10 : _GEN_9; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_11 = 8'hb == pc ? code_11 : _GEN_10; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_12 = 8'hc == pc ? code_12 : _GEN_11; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_13 = 8'hd == pc ? code_13 : _GEN_12; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_14 = 8'he == pc ? code_14 : _GEN_13; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_15 = 8'hf == pc ? code_15 : _GEN_14; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_16 = 8'h10 == pc ? code_16 : _GEN_15; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_17 = 8'h11 == pc ? code_17 : _GEN_16; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_18 = 8'h12 == pc ? code_18 : _GEN_17; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_19 = 8'h13 == pc ? code_19 : _GEN_18; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_20 = 8'h14 == pc ? code_20 : _GEN_19; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_21 = 8'h15 == pc ? code_21 : _GEN_20; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_22 = 8'h16 == pc ? code_22 : _GEN_21; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_23 = 8'h17 == pc ? code_23 : _GEN_22; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_24 = 8'h18 == pc ? code_24 : _GEN_23; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_25 = 8'h19 == pc ? code_25 : _GEN_24; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_26 = 8'h1a == pc ? code_26 : _GEN_25; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_27 = 8'h1b == pc ? code_27 : _GEN_26; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_28 = 8'h1c == pc ? code_28 : _GEN_27; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_29 = 8'h1d == pc ? code_29 : _GEN_28; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_30 = 8'h1e == pc ? code_30 : _GEN_29; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_31 = 8'h1f == pc ? code_31 : _GEN_30; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_32 = 8'h20 == pc ? code_32 : _GEN_31; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_33 = 8'h21 == pc ? code_33 : _GEN_32; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_34 = 8'h22 == pc ? code_34 : _GEN_33; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_35 = 8'h23 == pc ? code_35 : _GEN_34; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_36 = 8'h24 == pc ? code_36 : _GEN_35; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_37 = 8'h25 == pc ? code_37 : _GEN_36; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_38 = 8'h26 == pc ? code_38 : _GEN_37; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_39 = 8'h27 == pc ? code_39 : _GEN_38; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_40 = 8'h28 == pc ? code_40 : _GEN_39; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_41 = 8'h29 == pc ? code_41 : _GEN_40; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_42 = 8'h2a == pc ? code_42 : _GEN_41; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_43 = 8'h2b == pc ? code_43 : _GEN_42; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_44 = 8'h2c == pc ? code_44 : _GEN_43; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_45 = 8'h2d == pc ? code_45 : _GEN_44; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_46 = 8'h2e == pc ? code_46 : _GEN_45; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_47 = 8'h2f == pc ? code_47 : _GEN_46; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_48 = 8'h30 == pc ? code_48 : _GEN_47; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_49 = 8'h31 == pc ? code_49 : _GEN_48; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_50 = 8'h32 == pc ? code_50 : _GEN_49; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_51 = 8'h33 == pc ? code_51 : _GEN_50; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_52 = 8'h34 == pc ? code_52 : _GEN_51; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_53 = 8'h35 == pc ? code_53 : _GEN_52; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_54 = 8'h36 == pc ? code_54 : _GEN_53; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_55 = 8'h37 == pc ? code_55 : _GEN_54; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_56 = 8'h38 == pc ? code_56 : _GEN_55; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_57 = 8'h39 == pc ? code_57 : _GEN_56; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_58 = 8'h3a == pc ? code_58 : _GEN_57; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_59 = 8'h3b == pc ? code_59 : _GEN_58; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_60 = 8'h3c == pc ? code_60 : _GEN_59; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_61 = 8'h3d == pc ? code_61 : _GEN_60; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_62 = 8'h3e == pc ? code_62 : _GEN_61; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_63 = 8'h3f == pc ? code_63 : _GEN_62; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_64 = 8'h40 == pc ? code_64 : _GEN_63; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_65 = 8'h41 == pc ? code_65 : _GEN_64; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_66 = 8'h42 == pc ? code_66 : _GEN_65; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_67 = 8'h43 == pc ? code_67 : _GEN_66; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_68 = 8'h44 == pc ? code_68 : _GEN_67; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_69 = 8'h45 == pc ? code_69 : _GEN_68; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_70 = 8'h46 == pc ? code_70 : _GEN_69; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_71 = 8'h47 == pc ? code_71 : _GEN_70; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_72 = 8'h48 == pc ? code_72 : _GEN_71; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_73 = 8'h49 == pc ? code_73 : _GEN_72; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_74 = 8'h4a == pc ? code_74 : _GEN_73; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_75 = 8'h4b == pc ? code_75 : _GEN_74; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_76 = 8'h4c == pc ? code_76 : _GEN_75; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_77 = 8'h4d == pc ? code_77 : _GEN_76; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_78 = 8'h4e == pc ? code_78 : _GEN_77; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_79 = 8'h4f == pc ? code_79 : _GEN_78; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_80 = 8'h50 == pc ? code_80 : _GEN_79; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_81 = 8'h51 == pc ? code_81 : _GEN_80; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_82 = 8'h52 == pc ? code_82 : _GEN_81; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_83 = 8'h53 == pc ? code_83 : _GEN_82; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_84 = 8'h54 == pc ? code_84 : _GEN_83; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_85 = 8'h55 == pc ? code_85 : _GEN_84; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_86 = 8'h56 == pc ? code_86 : _GEN_85; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_87 = 8'h57 == pc ? code_87 : _GEN_86; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_88 = 8'h58 == pc ? code_88 : _GEN_87; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_89 = 8'h59 == pc ? code_89 : _GEN_88; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_90 = 8'h5a == pc ? code_90 : _GEN_89; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_91 = 8'h5b == pc ? code_91 : _GEN_90; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_92 = 8'h5c == pc ? code_92 : _GEN_91; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_93 = 8'h5d == pc ? code_93 : _GEN_92; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_94 = 8'h5e == pc ? code_94 : _GEN_93; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_95 = 8'h5f == pc ? code_95 : _GEN_94; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_96 = 8'h60 == pc ? code_96 : _GEN_95; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_97 = 8'h61 == pc ? code_97 : _GEN_96; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_98 = 8'h62 == pc ? code_98 : _GEN_97; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_99 = 8'h63 == pc ? code_99 : _GEN_98; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_100 = 8'h64 == pc ? code_100 : _GEN_99; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_101 = 8'h65 == pc ? code_101 : _GEN_100; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_102 = 8'h66 == pc ? code_102 : _GEN_101; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_103 = 8'h67 == pc ? code_103 : _GEN_102; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_104 = 8'h68 == pc ? code_104 : _GEN_103; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_105 = 8'h69 == pc ? code_105 : _GEN_104; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_106 = 8'h6a == pc ? code_106 : _GEN_105; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_107 = 8'h6b == pc ? code_107 : _GEN_106; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_108 = 8'h6c == pc ? code_108 : _GEN_107; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_109 = 8'h6d == pc ? code_109 : _GEN_108; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_110 = 8'h6e == pc ? code_110 : _GEN_109; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_111 = 8'h6f == pc ? code_111 : _GEN_110; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_112 = 8'h70 == pc ? code_112 : _GEN_111; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_113 = 8'h71 == pc ? code_113 : _GEN_112; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_114 = 8'h72 == pc ? code_114 : _GEN_113; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_115 = 8'h73 == pc ? code_115 : _GEN_114; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_116 = 8'h74 == pc ? code_116 : _GEN_115; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_117 = 8'h75 == pc ? code_117 : _GEN_116; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_118 = 8'h76 == pc ? code_118 : _GEN_117; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_119 = 8'h77 == pc ? code_119 : _GEN_118; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_120 = 8'h78 == pc ? code_120 : _GEN_119; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_121 = 8'h79 == pc ? code_121 : _GEN_120; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_122 = 8'h7a == pc ? code_122 : _GEN_121; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_123 = 8'h7b == pc ? code_123 : _GEN_122; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_124 = 8'h7c == pc ? code_124 : _GEN_123; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_125 = 8'h7d == pc ? code_125 : _GEN_124; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_126 = 8'h7e == pc ? code_126 : _GEN_125; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_127 = 8'h7f == pc ? code_127 : _GEN_126; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_128 = 8'h80 == pc ? code_128 : _GEN_127; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_129 = 8'h81 == pc ? code_129 : _GEN_128; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_130 = 8'h82 == pc ? code_130 : _GEN_129; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_131 = 8'h83 == pc ? code_131 : _GEN_130; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_132 = 8'h84 == pc ? code_132 : _GEN_131; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_133 = 8'h85 == pc ? code_133 : _GEN_132; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_134 = 8'h86 == pc ? code_134 : _GEN_133; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_135 = 8'h87 == pc ? code_135 : _GEN_134; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_136 = 8'h88 == pc ? code_136 : _GEN_135; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_137 = 8'h89 == pc ? code_137 : _GEN_136; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_138 = 8'h8a == pc ? code_138 : _GEN_137; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_139 = 8'h8b == pc ? code_139 : _GEN_138; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_140 = 8'h8c == pc ? code_140 : _GEN_139; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_141 = 8'h8d == pc ? code_141 : _GEN_140; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_142 = 8'h8e == pc ? code_142 : _GEN_141; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_143 = 8'h8f == pc ? code_143 : _GEN_142; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_144 = 8'h90 == pc ? code_144 : _GEN_143; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_145 = 8'h91 == pc ? code_145 : _GEN_144; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_146 = 8'h92 == pc ? code_146 : _GEN_145; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_147 = 8'h93 == pc ? code_147 : _GEN_146; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_148 = 8'h94 == pc ? code_148 : _GEN_147; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_149 = 8'h95 == pc ? code_149 : _GEN_148; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_150 = 8'h96 == pc ? code_150 : _GEN_149; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_151 = 8'h97 == pc ? code_151 : _GEN_150; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_152 = 8'h98 == pc ? code_152 : _GEN_151; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_153 = 8'h99 == pc ? code_153 : _GEN_152; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_154 = 8'h9a == pc ? code_154 : _GEN_153; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_155 = 8'h9b == pc ? code_155 : _GEN_154; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_156 = 8'h9c == pc ? code_156 : _GEN_155; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_157 = 8'h9d == pc ? code_157 : _GEN_156; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_158 = 8'h9e == pc ? code_158 : _GEN_157; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_159 = 8'h9f == pc ? code_159 : _GEN_158; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_160 = 8'ha0 == pc ? code_160 : _GEN_159; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_161 = 8'ha1 == pc ? code_161 : _GEN_160; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_162 = 8'ha2 == pc ? code_162 : _GEN_161; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_163 = 8'ha3 == pc ? code_163 : _GEN_162; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_164 = 8'ha4 == pc ? code_164 : _GEN_163; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_165 = 8'ha5 == pc ? code_165 : _GEN_164; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_166 = 8'ha6 == pc ? code_166 : _GEN_165; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_167 = 8'ha7 == pc ? code_167 : _GEN_166; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_168 = 8'ha8 == pc ? code_168 : _GEN_167; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_169 = 8'ha9 == pc ? code_169 : _GEN_168; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_170 = 8'haa == pc ? code_170 : _GEN_169; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_171 = 8'hab == pc ? code_171 : _GEN_170; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_172 = 8'hac == pc ? code_172 : _GEN_171; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_173 = 8'had == pc ? code_173 : _GEN_172; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_174 = 8'hae == pc ? code_174 : _GEN_173; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_175 = 8'haf == pc ? code_175 : _GEN_174; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_176 = 8'hb0 == pc ? code_176 : _GEN_175; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_177 = 8'hb1 == pc ? code_177 : _GEN_176; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_178 = 8'hb2 == pc ? code_178 : _GEN_177; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_179 = 8'hb3 == pc ? code_179 : _GEN_178; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_180 = 8'hb4 == pc ? code_180 : _GEN_179; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_181 = 8'hb5 == pc ? code_181 : _GEN_180; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_182 = 8'hb6 == pc ? code_182 : _GEN_181; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_183 = 8'hb7 == pc ? code_183 : _GEN_182; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_184 = 8'hb8 == pc ? code_184 : _GEN_183; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_185 = 8'hb9 == pc ? code_185 : _GEN_184; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_186 = 8'hba == pc ? code_186 : _GEN_185; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_187 = 8'hbb == pc ? code_187 : _GEN_186; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_188 = 8'hbc == pc ? code_188 : _GEN_187; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_189 = 8'hbd == pc ? code_189 : _GEN_188; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_190 = 8'hbe == pc ? code_190 : _GEN_189; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_191 = 8'hbf == pc ? code_191 : _GEN_190; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_192 = 8'hc0 == pc ? code_192 : _GEN_191; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_193 = 8'hc1 == pc ? code_193 : _GEN_192; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_194 = 8'hc2 == pc ? code_194 : _GEN_193; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_195 = 8'hc3 == pc ? code_195 : _GEN_194; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_196 = 8'hc4 == pc ? code_196 : _GEN_195; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_197 = 8'hc5 == pc ? code_197 : _GEN_196; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_198 = 8'hc6 == pc ? code_198 : _GEN_197; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_199 = 8'hc7 == pc ? code_199 : _GEN_198; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_200 = 8'hc8 == pc ? code_200 : _GEN_199; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_201 = 8'hc9 == pc ? code_201 : _GEN_200; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_202 = 8'hca == pc ? code_202 : _GEN_201; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_203 = 8'hcb == pc ? code_203 : _GEN_202; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_204 = 8'hcc == pc ? code_204 : _GEN_203; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_205 = 8'hcd == pc ? code_205 : _GEN_204; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_206 = 8'hce == pc ? code_206 : _GEN_205; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_207 = 8'hcf == pc ? code_207 : _GEN_206; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_208 = 8'hd0 == pc ? code_208 : _GEN_207; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_209 = 8'hd1 == pc ? code_209 : _GEN_208; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_210 = 8'hd2 == pc ? code_210 : _GEN_209; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_211 = 8'hd3 == pc ? code_211 : _GEN_210; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_212 = 8'hd4 == pc ? code_212 : _GEN_211; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_213 = 8'hd5 == pc ? code_213 : _GEN_212; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_214 = 8'hd6 == pc ? code_214 : _GEN_213; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_215 = 8'hd7 == pc ? code_215 : _GEN_214; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_216 = 8'hd8 == pc ? code_216 : _GEN_215; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_217 = 8'hd9 == pc ? code_217 : _GEN_216; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_218 = 8'hda == pc ? code_218 : _GEN_217; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_219 = 8'hdb == pc ? code_219 : _GEN_218; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_220 = 8'hdc == pc ? code_220 : _GEN_219; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_221 = 8'hdd == pc ? code_221 : _GEN_220; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_222 = 8'hde == pc ? code_222 : _GEN_221; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_223 = 8'hdf == pc ? code_223 : _GEN_222; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_224 = 8'he0 == pc ? code_224 : _GEN_223; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_225 = 8'he1 == pc ? code_225 : _GEN_224; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_226 = 8'he2 == pc ? code_226 : _GEN_225; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_227 = 8'he3 == pc ? code_227 : _GEN_226; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_228 = 8'he4 == pc ? code_228 : _GEN_227; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_229 = 8'he5 == pc ? code_229 : _GEN_228; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_230 = 8'he6 == pc ? code_230 : _GEN_229; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_231 = 8'he7 == pc ? code_231 : _GEN_230; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_232 = 8'he8 == pc ? code_232 : _GEN_231; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_233 = 8'he9 == pc ? code_233 : _GEN_232; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_234 = 8'hea == pc ? code_234 : _GEN_233; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_235 = 8'heb == pc ? code_235 : _GEN_234; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_236 = 8'hec == pc ? code_236 : _GEN_235; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_237 = 8'hed == pc ? code_237 : _GEN_236; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_238 = 8'hee == pc ? code_238 : _GEN_237; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_239 = 8'hef == pc ? code_239 : _GEN_238; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_240 = 8'hf0 == pc ? code_240 : _GEN_239; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_241 = 8'hf1 == pc ? code_241 : _GEN_240; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_242 = 8'hf2 == pc ? code_242 : _GEN_241; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_243 = 8'hf3 == pc ? code_243 : _GEN_242; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_244 = 8'hf4 == pc ? code_244 : _GEN_243; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_245 = 8'hf5 == pc ? code_245 : _GEN_244; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_246 = 8'hf6 == pc ? code_246 : _GEN_245; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_247 = 8'hf7 == pc ? code_247 : _GEN_246; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_248 = 8'hf8 == pc ? code_248 : _GEN_247; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_249 = 8'hf9 == pc ? code_249 : _GEN_248; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_250 = 8'hfa == pc ? code_250 : _GEN_249; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_251 = 8'hfb == pc ? code_251 : _GEN_250; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_252 = 8'hfc == pc ? code_252 : _GEN_251; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_253 = 8'hfd == pc ? code_253 : _GEN_252; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_254 = 8'hfe == pc ? code_254 : _GEN_253; // @[Risc.scala 27:{18,18}]
  wire [31:0] _GEN_255 = 8'hff == pc ? code_255 : _GEN_254; // @[Risc.scala 27:{18,18}]
  wire [7:0] op = _GEN_255[31:24]; // @[Risc.scala 27:18]
  wire [7:0] rci = _GEN_255[23:16]; // @[Risc.scala 28:18]
  wire [7:0] rai = _GEN_255[15:8]; // @[Risc.scala 29:18]
  wire [7:0] rbi = _GEN_255[7:0]; // @[Risc.scala 30:18]
  wire [31:0] ra = rai == 8'h0 ? 32'h0 : file_ra_MPORT_data; // @[Risc.scala 32:15]
  wire [31:0] rb = rbi == 8'h0 ? 32'h0 : file_rb_MPORT_data; // @[Risc.scala 33:15]
  wire [31:0] _rc_T_1 = ra + rb; // @[Risc.scala 46:29]
  wire [7:0] _rc_T_3 = rai + rbi; // @[Risc.scala 47:31]
  wire [7:0] _GEN_512 = 8'h1 == op ? _rc_T_3 : 8'h0; // @[Risc.scala 38:12 45:16 47:23]
  wire [31:0] _GEN_513 = 8'h33 == op ? _rc_T_1 : {{24'd0}, _GEN_512}; // @[Risc.scala 45:16 46:23]
  wire  _T_2 = rci == 8'hff; // @[Risc.scala 50:15]
  wire  _GEN_517 = rci == 8'hff ? 1'h0 : 1'h1; // @[Risc.scala 16:17 50:26 53:11]
  wire [31:0] _GEN_521 = io_boot ? 32'h0 : _GEN_513; // @[Risc.scala 38:12 42:25]
  wire [31:0] rc = io_isWr ? 32'h0 : _GEN_521; // @[Risc.scala 38:12 40:18]
  wire [7:0] _pc_T_1 = pc + 8'h1; // @[Risc.scala 55:14]
  wire [31:0] _GEN_522 = io_boot ? 32'h0 : rc; // @[Risc.scala 37:12 42:25 49:12]
  wire  _GEN_523 = io_boot ? 1'h0 : _T_2; // @[Risc.scala 36:12 42:25]
  wire  _GEN_526 = io_boot ? 1'h0 : _GEN_517; // @[Risc.scala 16:17 42:25]
  assign file_ra_MPORT_en = 1'h1;
  assign file_ra_MPORT_addr = _GEN_255[15:8];
  assign file_ra_MPORT_data = file[file_ra_MPORT_addr]; // @[Risc.scala 16:17]
  assign file_rb_MPORT_en = 1'h1;
  assign file_rb_MPORT_addr = _GEN_255[7:0];
  assign file_rb_MPORT_data = file[file_rb_MPORT_addr]; // @[Risc.scala 16:17]
  assign file_MPORT_data = io_isWr ? 32'h0 : _GEN_521;
  assign file_MPORT_addr = _GEN_255[23:16];
  assign file_MPORT_mask = 1'h1;
  assign file_MPORT_en = io_isWr ? 1'h0 : _GEN_526;
  assign io_valid = io_isWr ? 1'h0 : _GEN_523; // @[Risc.scala 36:12 40:18]
  assign io_out = io_isWr ? 32'h0 : _GEN_522; // @[Risc.scala 37:12 40:18]
  always @(posedge clock) begin
    if (file_MPORT_en & file_MPORT_mask) begin
      file[file_MPORT_addr] <= file_MPORT_data; // @[Risc.scala 16:17]
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_0 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h0 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_0 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_1 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h1 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_1 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_2 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h2 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_2 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_3 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h3 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_3 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_4 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h4 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_4 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_5 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h5 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_5 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_6 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h6 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_6 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_7 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h7 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_7 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_8 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h8 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_8 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_9 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h9 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_9 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_10 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'ha == io_wrAddr) begin // @[Risc.scala 41:21]
        code_10 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_11 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hb == io_wrAddr) begin // @[Risc.scala 41:21]
        code_11 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_12 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hc == io_wrAddr) begin // @[Risc.scala 41:21]
        code_12 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_13 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hd == io_wrAddr) begin // @[Risc.scala 41:21]
        code_13 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_14 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'he == io_wrAddr) begin // @[Risc.scala 41:21]
        code_14 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_15 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hf == io_wrAddr) begin // @[Risc.scala 41:21]
        code_15 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_16 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h10 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_16 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_17 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h11 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_17 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_18 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h12 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_18 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_19 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h13 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_19 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_20 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h14 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_20 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_21 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h15 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_21 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_22 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h16 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_22 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_23 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h17 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_23 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_24 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h18 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_24 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_25 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h19 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_25 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_26 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h1a == io_wrAddr) begin // @[Risc.scala 41:21]
        code_26 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_27 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h1b == io_wrAddr) begin // @[Risc.scala 41:21]
        code_27 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_28 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h1c == io_wrAddr) begin // @[Risc.scala 41:21]
        code_28 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_29 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h1d == io_wrAddr) begin // @[Risc.scala 41:21]
        code_29 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_30 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h1e == io_wrAddr) begin // @[Risc.scala 41:21]
        code_30 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_31 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h1f == io_wrAddr) begin // @[Risc.scala 41:21]
        code_31 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_32 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h20 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_32 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_33 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h21 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_33 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_34 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h22 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_34 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_35 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h23 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_35 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_36 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h24 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_36 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_37 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h25 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_37 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_38 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h26 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_38 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_39 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h27 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_39 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_40 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h28 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_40 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_41 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h29 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_41 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_42 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h2a == io_wrAddr) begin // @[Risc.scala 41:21]
        code_42 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_43 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h2b == io_wrAddr) begin // @[Risc.scala 41:21]
        code_43 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_44 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h2c == io_wrAddr) begin // @[Risc.scala 41:21]
        code_44 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_45 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h2d == io_wrAddr) begin // @[Risc.scala 41:21]
        code_45 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_46 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h2e == io_wrAddr) begin // @[Risc.scala 41:21]
        code_46 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_47 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h2f == io_wrAddr) begin // @[Risc.scala 41:21]
        code_47 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_48 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h30 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_48 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_49 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h31 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_49 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_50 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h32 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_50 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_51 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h33 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_51 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_52 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h34 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_52 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_53 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h35 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_53 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_54 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h36 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_54 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_55 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h37 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_55 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_56 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h38 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_56 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_57 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h39 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_57 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_58 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h3a == io_wrAddr) begin // @[Risc.scala 41:21]
        code_58 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_59 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h3b == io_wrAddr) begin // @[Risc.scala 41:21]
        code_59 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_60 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h3c == io_wrAddr) begin // @[Risc.scala 41:21]
        code_60 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_61 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h3d == io_wrAddr) begin // @[Risc.scala 41:21]
        code_61 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_62 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h3e == io_wrAddr) begin // @[Risc.scala 41:21]
        code_62 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_63 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h3f == io_wrAddr) begin // @[Risc.scala 41:21]
        code_63 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_64 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h40 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_64 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_65 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h41 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_65 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_66 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h42 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_66 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_67 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h43 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_67 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_68 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h44 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_68 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_69 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h45 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_69 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_70 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h46 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_70 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_71 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h47 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_71 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_72 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h48 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_72 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_73 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h49 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_73 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_74 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h4a == io_wrAddr) begin // @[Risc.scala 41:21]
        code_74 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_75 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h4b == io_wrAddr) begin // @[Risc.scala 41:21]
        code_75 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_76 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h4c == io_wrAddr) begin // @[Risc.scala 41:21]
        code_76 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_77 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h4d == io_wrAddr) begin // @[Risc.scala 41:21]
        code_77 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_78 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h4e == io_wrAddr) begin // @[Risc.scala 41:21]
        code_78 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_79 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h4f == io_wrAddr) begin // @[Risc.scala 41:21]
        code_79 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_80 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h50 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_80 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_81 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h51 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_81 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_82 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h52 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_82 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_83 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h53 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_83 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_84 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h54 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_84 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_85 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h55 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_85 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_86 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h56 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_86 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_87 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h57 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_87 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_88 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h58 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_88 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_89 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h59 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_89 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_90 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h5a == io_wrAddr) begin // @[Risc.scala 41:21]
        code_90 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_91 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h5b == io_wrAddr) begin // @[Risc.scala 41:21]
        code_91 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_92 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h5c == io_wrAddr) begin // @[Risc.scala 41:21]
        code_92 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_93 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h5d == io_wrAddr) begin // @[Risc.scala 41:21]
        code_93 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_94 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h5e == io_wrAddr) begin // @[Risc.scala 41:21]
        code_94 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_95 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h5f == io_wrAddr) begin // @[Risc.scala 41:21]
        code_95 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_96 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h60 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_96 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_97 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h61 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_97 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_98 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h62 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_98 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_99 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h63 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_99 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_100 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h64 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_100 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_101 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h65 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_101 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_102 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h66 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_102 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_103 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h67 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_103 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_104 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h68 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_104 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_105 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h69 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_105 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_106 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h6a == io_wrAddr) begin // @[Risc.scala 41:21]
        code_106 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_107 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h6b == io_wrAddr) begin // @[Risc.scala 41:21]
        code_107 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_108 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h6c == io_wrAddr) begin // @[Risc.scala 41:21]
        code_108 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_109 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h6d == io_wrAddr) begin // @[Risc.scala 41:21]
        code_109 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_110 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h6e == io_wrAddr) begin // @[Risc.scala 41:21]
        code_110 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_111 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h6f == io_wrAddr) begin // @[Risc.scala 41:21]
        code_111 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_112 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h70 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_112 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_113 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h71 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_113 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_114 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h72 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_114 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_115 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h73 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_115 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_116 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h74 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_116 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_117 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h75 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_117 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_118 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h76 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_118 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_119 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h77 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_119 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_120 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h78 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_120 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_121 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h79 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_121 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_122 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h7a == io_wrAddr) begin // @[Risc.scala 41:21]
        code_122 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_123 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h7b == io_wrAddr) begin // @[Risc.scala 41:21]
        code_123 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_124 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h7c == io_wrAddr) begin // @[Risc.scala 41:21]
        code_124 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_125 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h7d == io_wrAddr) begin // @[Risc.scala 41:21]
        code_125 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_126 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h7e == io_wrAddr) begin // @[Risc.scala 41:21]
        code_126 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_127 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h7f == io_wrAddr) begin // @[Risc.scala 41:21]
        code_127 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_128 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h80 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_128 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_129 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h81 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_129 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_130 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h82 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_130 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_131 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h83 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_131 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_132 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h84 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_132 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_133 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h85 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_133 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_134 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h86 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_134 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_135 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h87 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_135 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_136 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h88 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_136 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_137 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h89 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_137 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_138 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h8a == io_wrAddr) begin // @[Risc.scala 41:21]
        code_138 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_139 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h8b == io_wrAddr) begin // @[Risc.scala 41:21]
        code_139 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_140 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h8c == io_wrAddr) begin // @[Risc.scala 41:21]
        code_140 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_141 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h8d == io_wrAddr) begin // @[Risc.scala 41:21]
        code_141 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_142 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h8e == io_wrAddr) begin // @[Risc.scala 41:21]
        code_142 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_143 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h8f == io_wrAddr) begin // @[Risc.scala 41:21]
        code_143 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_144 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h90 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_144 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_145 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h91 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_145 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_146 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h92 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_146 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_147 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h93 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_147 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_148 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h94 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_148 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_149 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h95 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_149 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_150 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h96 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_150 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_151 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h97 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_151 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_152 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h98 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_152 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_153 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h99 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_153 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_154 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h9a == io_wrAddr) begin // @[Risc.scala 41:21]
        code_154 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_155 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h9b == io_wrAddr) begin // @[Risc.scala 41:21]
        code_155 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_156 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h9c == io_wrAddr) begin // @[Risc.scala 41:21]
        code_156 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_157 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h9d == io_wrAddr) begin // @[Risc.scala 41:21]
        code_157 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_158 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h9e == io_wrAddr) begin // @[Risc.scala 41:21]
        code_158 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_159 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'h9f == io_wrAddr) begin // @[Risc.scala 41:21]
        code_159 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_160 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'ha0 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_160 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_161 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'ha1 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_161 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_162 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'ha2 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_162 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_163 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'ha3 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_163 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_164 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'ha4 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_164 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_165 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'ha5 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_165 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_166 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'ha6 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_166 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_167 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'ha7 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_167 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_168 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'ha8 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_168 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_169 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'ha9 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_169 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_170 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'haa == io_wrAddr) begin // @[Risc.scala 41:21]
        code_170 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_171 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hab == io_wrAddr) begin // @[Risc.scala 41:21]
        code_171 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_172 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hac == io_wrAddr) begin // @[Risc.scala 41:21]
        code_172 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_173 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'had == io_wrAddr) begin // @[Risc.scala 41:21]
        code_173 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_174 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hae == io_wrAddr) begin // @[Risc.scala 41:21]
        code_174 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_175 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'haf == io_wrAddr) begin // @[Risc.scala 41:21]
        code_175 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_176 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hb0 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_176 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_177 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hb1 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_177 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_178 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hb2 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_178 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_179 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hb3 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_179 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_180 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hb4 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_180 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_181 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hb5 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_181 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_182 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hb6 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_182 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_183 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hb7 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_183 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_184 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hb8 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_184 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_185 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hb9 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_185 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_186 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hba == io_wrAddr) begin // @[Risc.scala 41:21]
        code_186 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_187 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hbb == io_wrAddr) begin // @[Risc.scala 41:21]
        code_187 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_188 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hbc == io_wrAddr) begin // @[Risc.scala 41:21]
        code_188 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_189 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hbd == io_wrAddr) begin // @[Risc.scala 41:21]
        code_189 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_190 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hbe == io_wrAddr) begin // @[Risc.scala 41:21]
        code_190 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_191 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hbf == io_wrAddr) begin // @[Risc.scala 41:21]
        code_191 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_192 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hc0 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_192 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_193 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hc1 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_193 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_194 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hc2 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_194 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_195 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hc3 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_195 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_196 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hc4 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_196 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_197 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hc5 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_197 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_198 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hc6 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_198 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_199 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hc7 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_199 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_200 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hc8 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_200 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_201 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hc9 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_201 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_202 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hca == io_wrAddr) begin // @[Risc.scala 41:21]
        code_202 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_203 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hcb == io_wrAddr) begin // @[Risc.scala 41:21]
        code_203 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_204 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hcc == io_wrAddr) begin // @[Risc.scala 41:21]
        code_204 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_205 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hcd == io_wrAddr) begin // @[Risc.scala 41:21]
        code_205 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_206 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hce == io_wrAddr) begin // @[Risc.scala 41:21]
        code_206 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_207 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hcf == io_wrAddr) begin // @[Risc.scala 41:21]
        code_207 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_208 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hd0 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_208 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_209 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hd1 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_209 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_210 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hd2 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_210 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_211 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hd3 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_211 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_212 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hd4 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_212 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_213 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hd5 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_213 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_214 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hd6 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_214 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_215 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hd7 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_215 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_216 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hd8 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_216 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_217 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hd9 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_217 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_218 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hda == io_wrAddr) begin // @[Risc.scala 41:21]
        code_218 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_219 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hdb == io_wrAddr) begin // @[Risc.scala 41:21]
        code_219 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_220 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hdc == io_wrAddr) begin // @[Risc.scala 41:21]
        code_220 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_221 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hdd == io_wrAddr) begin // @[Risc.scala 41:21]
        code_221 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_222 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hde == io_wrAddr) begin // @[Risc.scala 41:21]
        code_222 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_223 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hdf == io_wrAddr) begin // @[Risc.scala 41:21]
        code_223 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_224 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'he0 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_224 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_225 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'he1 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_225 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_226 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'he2 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_226 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_227 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'he3 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_227 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_228 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'he4 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_228 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_229 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'he5 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_229 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_230 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'he6 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_230 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_231 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'he7 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_231 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_232 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'he8 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_232 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_233 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'he9 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_233 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_234 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hea == io_wrAddr) begin // @[Risc.scala 41:21]
        code_234 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_235 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'heb == io_wrAddr) begin // @[Risc.scala 41:21]
        code_235 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_236 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hec == io_wrAddr) begin // @[Risc.scala 41:21]
        code_236 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_237 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hed == io_wrAddr) begin // @[Risc.scala 41:21]
        code_237 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_238 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hee == io_wrAddr) begin // @[Risc.scala 41:21]
        code_238 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_239 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hef == io_wrAddr) begin // @[Risc.scala 41:21]
        code_239 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_240 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hf0 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_240 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_241 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hf1 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_241 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_242 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hf2 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_242 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_243 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hf3 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_243 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_244 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hf4 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_244 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_245 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hf5 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_245 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_246 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hf6 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_246 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_247 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hf7 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_247 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_248 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hf8 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_248 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_249 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hf9 == io_wrAddr) begin // @[Risc.scala 41:21]
        code_249 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_250 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hfa == io_wrAddr) begin // @[Risc.scala 41:21]
        code_250 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_251 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hfb == io_wrAddr) begin // @[Risc.scala 41:21]
        code_251 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_252 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hfc == io_wrAddr) begin // @[Risc.scala 41:21]
        code_252 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_253 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hfd == io_wrAddr) begin // @[Risc.scala 41:21]
        code_253 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_254 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hfe == io_wrAddr) begin // @[Risc.scala 41:21]
        code_254 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 19:21]
      code_255 <= 32'h0; // @[Risc.scala 19:21]
    end else if (io_isWr) begin // @[Risc.scala 40:18]
      if (8'hff == io_wrAddr) begin // @[Risc.scala 41:21]
        code_255 <= io_wrData; // @[Risc.scala 41:21]
      end
    end
    if (reset) begin // @[Risc.scala 21:21]
      pc <= 8'h0; // @[Risc.scala 21:21]
    end else if (!(io_isWr)) begin // @[Risc.scala 40:18]
      if (io_boot) begin // @[Risc.scala 42:25]
        pc <= 8'h0; // @[Risc.scala 43:8]
      end else begin
        pc <= _pc_T_1; // @[Risc.scala 55:8]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    file[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  code_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  code_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  code_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  code_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  code_4 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  code_5 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  code_6 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  code_7 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  code_8 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  code_9 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  code_10 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  code_11 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  code_12 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  code_13 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  code_14 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  code_15 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  code_16 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  code_17 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  code_18 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  code_19 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  code_20 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  code_21 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  code_22 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  code_23 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  code_24 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  code_25 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  code_26 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  code_27 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  code_28 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  code_29 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  code_30 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  code_31 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  code_32 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  code_33 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  code_34 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  code_35 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  code_36 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  code_37 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  code_38 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  code_39 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  code_40 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  code_41 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  code_42 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  code_43 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  code_44 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  code_45 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  code_46 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  code_47 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  code_48 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  code_49 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  code_50 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  code_51 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  code_52 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  code_53 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  code_54 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  code_55 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  code_56 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  code_57 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  code_58 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  code_59 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  code_60 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  code_61 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  code_62 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  code_63 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  code_64 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  code_65 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  code_66 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  code_67 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  code_68 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  code_69 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  code_70 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  code_71 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  code_72 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  code_73 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  code_74 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  code_75 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  code_76 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  code_77 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  code_78 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  code_79 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  code_80 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  code_81 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  code_82 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  code_83 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  code_84 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  code_85 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  code_86 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  code_87 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  code_88 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  code_89 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  code_90 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  code_91 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  code_92 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  code_93 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  code_94 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  code_95 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  code_96 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  code_97 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  code_98 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  code_99 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  code_100 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  code_101 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  code_102 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  code_103 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  code_104 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  code_105 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  code_106 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  code_107 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  code_108 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  code_109 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  code_110 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  code_111 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  code_112 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  code_113 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  code_114 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  code_115 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  code_116 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  code_117 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  code_118 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  code_119 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  code_120 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  code_121 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  code_122 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  code_123 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  code_124 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  code_125 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  code_126 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  code_127 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  code_128 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  code_129 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  code_130 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  code_131 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  code_132 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  code_133 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  code_134 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  code_135 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  code_136 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  code_137 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  code_138 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  code_139 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  code_140 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  code_141 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  code_142 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  code_143 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  code_144 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  code_145 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  code_146 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  code_147 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  code_148 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  code_149 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  code_150 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  code_151 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  code_152 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  code_153 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  code_154 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  code_155 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  code_156 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  code_157 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  code_158 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  code_159 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  code_160 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  code_161 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  code_162 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  code_163 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  code_164 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  code_165 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  code_166 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  code_167 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  code_168 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  code_169 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  code_170 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  code_171 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  code_172 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  code_173 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  code_174 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  code_175 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  code_176 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  code_177 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  code_178 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  code_179 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  code_180 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  code_181 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  code_182 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  code_183 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  code_184 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  code_185 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  code_186 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  code_187 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  code_188 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  code_189 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  code_190 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  code_191 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  code_192 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  code_193 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  code_194 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  code_195 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  code_196 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  code_197 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  code_198 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  code_199 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  code_200 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  code_201 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  code_202 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  code_203 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  code_204 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  code_205 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  code_206 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  code_207 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  code_208 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  code_209 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  code_210 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  code_211 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  code_212 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  code_213 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  code_214 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  code_215 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  code_216 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  code_217 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  code_218 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  code_219 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  code_220 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  code_221 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  code_222 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  code_223 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  code_224 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  code_225 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  code_226 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  code_227 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  code_228 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  code_229 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  code_230 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  code_231 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  code_232 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  code_233 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  code_234 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  code_235 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  code_236 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  code_237 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  code_238 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  code_239 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  code_240 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  code_241 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  code_242 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  code_243 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  code_244 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  code_245 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  code_246 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  code_247 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  code_248 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  code_249 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  code_250 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  code_251 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  code_252 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  code_253 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  code_254 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  code_255 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  pc = _RAND_257[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
