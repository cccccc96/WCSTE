module RISCVCPUv2(
  input         clock,
  input         reset,
  input  [4:0]  io_rvfi_rs1_addr_in,
  input  [4:0]  io_rvfi_rs2_addr_in,
  input  [63:0] io_rvfi_rs1_rdata_in,
  input  [63:0] io_rvfi_rs2_rdata_in,
  input         io_rvfi_rst,
  input  [31:0] io_rvfi_insn_in_0,
  input  [31:0] io_rvfi_insn_in_1,
  input  [31:0] io_rvfi_insn_in_2,
  input  [31:0] io_rvfi_insn_in_3,
  input  [9:0]  io_rvfi_mem_addr_in_0,
  input  [9:0]  io_rvfi_mem_addr_in_1,
  input  [31:0] io_rvfi_mem_data_in_0,
  input  [31:0] io_rvfi_mem_data_in_1,
  output        io_rvfi_valid,
  output [31:0] io_rvfi_insn,
  output [63:0] io_rvfi_pc_rdata,
  output [63:0] io_rvfi_pc_wdata,
  output [4:0]  io_rvfi_rs1_addr,
  output [4:0]  io_rvfi_rs2_addr,
  output [63:0] io_rvfi_rs1_rdata,
  output [63:0] io_rvfi_rs2_rdata,
  output [4:0]  io_rvfi_rd_addr,
  output [63:0] io_rvfi_rd_wdata,
  output [31:0] io_rvfi_mem_addr,
  output [63:0] io_rvfi_mem_rdata,
  output [63:0] io_rvfi_mem_wdata,
  output [63:0] io_rvfi_regs_0,
  output [63:0] io_rvfi_regs_1,
  output [63:0] io_rvfi_regs_2,
  output [63:0] io_rvfi_regs_3,
  output [63:0] io_rvfi_regs_4,
  output [63:0] io_rvfi_regs_5,
  output [63:0] io_rvfi_regs_6,
  output [63:0] io_rvfi_regs_7,
  output [63:0] io_rvfi_regs_8,
  output [63:0] io_rvfi_regs_9,
  output [63:0] io_rvfi_regs_10,
  output [63:0] io_rvfi_regs_11,
  output [63:0] io_rvfi_regs_12,
  output [63:0] io_rvfi_regs_13,
  output [63:0] io_rvfi_regs_14,
  output [63:0] io_rvfi_regs_15,
  output [63:0] io_rvfi_regs_16,
  output [63:0] io_rvfi_regs_17,
  output [63:0] io_rvfi_regs_18,
  output [63:0] io_rvfi_regs_19,
  output [63:0] io_rvfi_regs_20,
  output [63:0] io_rvfi_regs_21,
  output [63:0] io_rvfi_regs_22,
  output [63:0] io_rvfi_regs_23,
  output [63:0] io_rvfi_regs_24,
  output [63:0] io_rvfi_regs_25,
  output [63:0] io_rvfi_regs_26,
  output [63:0] io_rvfi_regs_27,
  output [63:0] io_rvfi_regs_28,
  output [63:0] io_rvfi_regs_29,
  output [63:0] io_rvfi_regs_30,
  output [63:0] io_rvfi_regs_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [63:0] _RAND_1070;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] PC; // @[CPU.scala 48:19]
  reg [63:0] Regs_0; // @[CPU.scala 49:17]
  reg [63:0] Regs_1; // @[CPU.scala 49:17]
  reg [63:0] Regs_2; // @[CPU.scala 49:17]
  reg [63:0] Regs_3; // @[CPU.scala 49:17]
  reg [63:0] Regs_4; // @[CPU.scala 49:17]
  reg [63:0] Regs_5; // @[CPU.scala 49:17]
  reg [63:0] Regs_6; // @[CPU.scala 49:17]
  reg [63:0] Regs_7; // @[CPU.scala 49:17]
  reg [63:0] Regs_8; // @[CPU.scala 49:17]
  reg [63:0] Regs_9; // @[CPU.scala 49:17]
  reg [63:0] Regs_10; // @[CPU.scala 49:17]
  reg [63:0] Regs_11; // @[CPU.scala 49:17]
  reg [63:0] Regs_12; // @[CPU.scala 49:17]
  reg [63:0] Regs_13; // @[CPU.scala 49:17]
  reg [63:0] Regs_14; // @[CPU.scala 49:17]
  reg [63:0] Regs_15; // @[CPU.scala 49:17]
  reg [63:0] Regs_16; // @[CPU.scala 49:17]
  reg [63:0] Regs_17; // @[CPU.scala 49:17]
  reg [63:0] Regs_18; // @[CPU.scala 49:17]
  reg [63:0] Regs_19; // @[CPU.scala 49:17]
  reg [63:0] Regs_20; // @[CPU.scala 49:17]
  reg [63:0] Regs_21; // @[CPU.scala 49:17]
  reg [63:0] Regs_22; // @[CPU.scala 49:17]
  reg [63:0] Regs_23; // @[CPU.scala 49:17]
  reg [63:0] Regs_24; // @[CPU.scala 49:17]
  reg [63:0] Regs_25; // @[CPU.scala 49:17]
  reg [63:0] Regs_26; // @[CPU.scala 49:17]
  reg [63:0] Regs_27; // @[CPU.scala 49:17]
  reg [63:0] Regs_28; // @[CPU.scala 49:17]
  reg [63:0] Regs_29; // @[CPU.scala 49:17]
  reg [63:0] Regs_30; // @[CPU.scala 49:17]
  reg [63:0] Regs_31; // @[CPU.scala 49:17]
  reg [63:0] IDEXA; // @[CPU.scala 50:58]
  reg [63:0] IDEXB; // @[CPU.scala 50:58]
  reg [63:0] EXMEMB; // @[CPU.scala 50:58]
  reg [63:0] EXMEMALUOut; // @[CPU.scala 50:58]
  reg [63:0] MEMWBValue; // @[CPU.scala 50:58]
  reg [31:0] DMemory_0; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1; // @[CPU.scala 52:20]
  reg [31:0] DMemory_2; // @[CPU.scala 52:20]
  reg [31:0] DMemory_3; // @[CPU.scala 52:20]
  reg [31:0] DMemory_4; // @[CPU.scala 52:20]
  reg [31:0] DMemory_5; // @[CPU.scala 52:20]
  reg [31:0] DMemory_6; // @[CPU.scala 52:20]
  reg [31:0] DMemory_7; // @[CPU.scala 52:20]
  reg [31:0] DMemory_8; // @[CPU.scala 52:20]
  reg [31:0] DMemory_9; // @[CPU.scala 52:20]
  reg [31:0] DMemory_10; // @[CPU.scala 52:20]
  reg [31:0] DMemory_11; // @[CPU.scala 52:20]
  reg [31:0] DMemory_12; // @[CPU.scala 52:20]
  reg [31:0] DMemory_13; // @[CPU.scala 52:20]
  reg [31:0] DMemory_14; // @[CPU.scala 52:20]
  reg [31:0] DMemory_15; // @[CPU.scala 52:20]
  reg [31:0] DMemory_16; // @[CPU.scala 52:20]
  reg [31:0] DMemory_17; // @[CPU.scala 52:20]
  reg [31:0] DMemory_18; // @[CPU.scala 52:20]
  reg [31:0] DMemory_19; // @[CPU.scala 52:20]
  reg [31:0] DMemory_20; // @[CPU.scala 52:20]
  reg [31:0] DMemory_21; // @[CPU.scala 52:20]
  reg [31:0] DMemory_22; // @[CPU.scala 52:20]
  reg [31:0] DMemory_23; // @[CPU.scala 52:20]
  reg [31:0] DMemory_24; // @[CPU.scala 52:20]
  reg [31:0] DMemory_25; // @[CPU.scala 52:20]
  reg [31:0] DMemory_26; // @[CPU.scala 52:20]
  reg [31:0] DMemory_27; // @[CPU.scala 52:20]
  reg [31:0] DMemory_28; // @[CPU.scala 52:20]
  reg [31:0] DMemory_29; // @[CPU.scala 52:20]
  reg [31:0] DMemory_30; // @[CPU.scala 52:20]
  reg [31:0] DMemory_31; // @[CPU.scala 52:20]
  reg [31:0] DMemory_32; // @[CPU.scala 52:20]
  reg [31:0] DMemory_33; // @[CPU.scala 52:20]
  reg [31:0] DMemory_34; // @[CPU.scala 52:20]
  reg [31:0] DMemory_35; // @[CPU.scala 52:20]
  reg [31:0] DMemory_36; // @[CPU.scala 52:20]
  reg [31:0] DMemory_37; // @[CPU.scala 52:20]
  reg [31:0] DMemory_38; // @[CPU.scala 52:20]
  reg [31:0] DMemory_39; // @[CPU.scala 52:20]
  reg [31:0] DMemory_40; // @[CPU.scala 52:20]
  reg [31:0] DMemory_41; // @[CPU.scala 52:20]
  reg [31:0] DMemory_42; // @[CPU.scala 52:20]
  reg [31:0] DMemory_43; // @[CPU.scala 52:20]
  reg [31:0] DMemory_44; // @[CPU.scala 52:20]
  reg [31:0] DMemory_45; // @[CPU.scala 52:20]
  reg [31:0] DMemory_46; // @[CPU.scala 52:20]
  reg [31:0] DMemory_47; // @[CPU.scala 52:20]
  reg [31:0] DMemory_48; // @[CPU.scala 52:20]
  reg [31:0] DMemory_49; // @[CPU.scala 52:20]
  reg [31:0] DMemory_50; // @[CPU.scala 52:20]
  reg [31:0] DMemory_51; // @[CPU.scala 52:20]
  reg [31:0] DMemory_52; // @[CPU.scala 52:20]
  reg [31:0] DMemory_53; // @[CPU.scala 52:20]
  reg [31:0] DMemory_54; // @[CPU.scala 52:20]
  reg [31:0] DMemory_55; // @[CPU.scala 52:20]
  reg [31:0] DMemory_56; // @[CPU.scala 52:20]
  reg [31:0] DMemory_57; // @[CPU.scala 52:20]
  reg [31:0] DMemory_58; // @[CPU.scala 52:20]
  reg [31:0] DMemory_59; // @[CPU.scala 52:20]
  reg [31:0] DMemory_60; // @[CPU.scala 52:20]
  reg [31:0] DMemory_61; // @[CPU.scala 52:20]
  reg [31:0] DMemory_62; // @[CPU.scala 52:20]
  reg [31:0] DMemory_63; // @[CPU.scala 52:20]
  reg [31:0] DMemory_64; // @[CPU.scala 52:20]
  reg [31:0] DMemory_65; // @[CPU.scala 52:20]
  reg [31:0] DMemory_66; // @[CPU.scala 52:20]
  reg [31:0] DMemory_67; // @[CPU.scala 52:20]
  reg [31:0] DMemory_68; // @[CPU.scala 52:20]
  reg [31:0] DMemory_69; // @[CPU.scala 52:20]
  reg [31:0] DMemory_70; // @[CPU.scala 52:20]
  reg [31:0] DMemory_71; // @[CPU.scala 52:20]
  reg [31:0] DMemory_72; // @[CPU.scala 52:20]
  reg [31:0] DMemory_73; // @[CPU.scala 52:20]
  reg [31:0] DMemory_74; // @[CPU.scala 52:20]
  reg [31:0] DMemory_75; // @[CPU.scala 52:20]
  reg [31:0] DMemory_76; // @[CPU.scala 52:20]
  reg [31:0] DMemory_77; // @[CPU.scala 52:20]
  reg [31:0] DMemory_78; // @[CPU.scala 52:20]
  reg [31:0] DMemory_79; // @[CPU.scala 52:20]
  reg [31:0] DMemory_80; // @[CPU.scala 52:20]
  reg [31:0] DMemory_81; // @[CPU.scala 52:20]
  reg [31:0] DMemory_82; // @[CPU.scala 52:20]
  reg [31:0] DMemory_83; // @[CPU.scala 52:20]
  reg [31:0] DMemory_84; // @[CPU.scala 52:20]
  reg [31:0] DMemory_85; // @[CPU.scala 52:20]
  reg [31:0] DMemory_86; // @[CPU.scala 52:20]
  reg [31:0] DMemory_87; // @[CPU.scala 52:20]
  reg [31:0] DMemory_88; // @[CPU.scala 52:20]
  reg [31:0] DMemory_89; // @[CPU.scala 52:20]
  reg [31:0] DMemory_90; // @[CPU.scala 52:20]
  reg [31:0] DMemory_91; // @[CPU.scala 52:20]
  reg [31:0] DMemory_92; // @[CPU.scala 52:20]
  reg [31:0] DMemory_93; // @[CPU.scala 52:20]
  reg [31:0] DMemory_94; // @[CPU.scala 52:20]
  reg [31:0] DMemory_95; // @[CPU.scala 52:20]
  reg [31:0] DMemory_96; // @[CPU.scala 52:20]
  reg [31:0] DMemory_97; // @[CPU.scala 52:20]
  reg [31:0] DMemory_98; // @[CPU.scala 52:20]
  reg [31:0] DMemory_99; // @[CPU.scala 52:20]
  reg [31:0] DMemory_100; // @[CPU.scala 52:20]
  reg [31:0] DMemory_101; // @[CPU.scala 52:20]
  reg [31:0] DMemory_102; // @[CPU.scala 52:20]
  reg [31:0] DMemory_103; // @[CPU.scala 52:20]
  reg [31:0] DMemory_104; // @[CPU.scala 52:20]
  reg [31:0] DMemory_105; // @[CPU.scala 52:20]
  reg [31:0] DMemory_106; // @[CPU.scala 52:20]
  reg [31:0] DMemory_107; // @[CPU.scala 52:20]
  reg [31:0] DMemory_108; // @[CPU.scala 52:20]
  reg [31:0] DMemory_109; // @[CPU.scala 52:20]
  reg [31:0] DMemory_110; // @[CPU.scala 52:20]
  reg [31:0] DMemory_111; // @[CPU.scala 52:20]
  reg [31:0] DMemory_112; // @[CPU.scala 52:20]
  reg [31:0] DMemory_113; // @[CPU.scala 52:20]
  reg [31:0] DMemory_114; // @[CPU.scala 52:20]
  reg [31:0] DMemory_115; // @[CPU.scala 52:20]
  reg [31:0] DMemory_116; // @[CPU.scala 52:20]
  reg [31:0] DMemory_117; // @[CPU.scala 52:20]
  reg [31:0] DMemory_118; // @[CPU.scala 52:20]
  reg [31:0] DMemory_119; // @[CPU.scala 52:20]
  reg [31:0] DMemory_120; // @[CPU.scala 52:20]
  reg [31:0] DMemory_121; // @[CPU.scala 52:20]
  reg [31:0] DMemory_122; // @[CPU.scala 52:20]
  reg [31:0] DMemory_123; // @[CPU.scala 52:20]
  reg [31:0] DMemory_124; // @[CPU.scala 52:20]
  reg [31:0] DMemory_125; // @[CPU.scala 52:20]
  reg [31:0] DMemory_126; // @[CPU.scala 52:20]
  reg [31:0] DMemory_127; // @[CPU.scala 52:20]
  reg [31:0] DMemory_128; // @[CPU.scala 52:20]
  reg [31:0] DMemory_129; // @[CPU.scala 52:20]
  reg [31:0] DMemory_130; // @[CPU.scala 52:20]
  reg [31:0] DMemory_131; // @[CPU.scala 52:20]
  reg [31:0] DMemory_132; // @[CPU.scala 52:20]
  reg [31:0] DMemory_133; // @[CPU.scala 52:20]
  reg [31:0] DMemory_134; // @[CPU.scala 52:20]
  reg [31:0] DMemory_135; // @[CPU.scala 52:20]
  reg [31:0] DMemory_136; // @[CPU.scala 52:20]
  reg [31:0] DMemory_137; // @[CPU.scala 52:20]
  reg [31:0] DMemory_138; // @[CPU.scala 52:20]
  reg [31:0] DMemory_139; // @[CPU.scala 52:20]
  reg [31:0] DMemory_140; // @[CPU.scala 52:20]
  reg [31:0] DMemory_141; // @[CPU.scala 52:20]
  reg [31:0] DMemory_142; // @[CPU.scala 52:20]
  reg [31:0] DMemory_143; // @[CPU.scala 52:20]
  reg [31:0] DMemory_144; // @[CPU.scala 52:20]
  reg [31:0] DMemory_145; // @[CPU.scala 52:20]
  reg [31:0] DMemory_146; // @[CPU.scala 52:20]
  reg [31:0] DMemory_147; // @[CPU.scala 52:20]
  reg [31:0] DMemory_148; // @[CPU.scala 52:20]
  reg [31:0] DMemory_149; // @[CPU.scala 52:20]
  reg [31:0] DMemory_150; // @[CPU.scala 52:20]
  reg [31:0] DMemory_151; // @[CPU.scala 52:20]
  reg [31:0] DMemory_152; // @[CPU.scala 52:20]
  reg [31:0] DMemory_153; // @[CPU.scala 52:20]
  reg [31:0] DMemory_154; // @[CPU.scala 52:20]
  reg [31:0] DMemory_155; // @[CPU.scala 52:20]
  reg [31:0] DMemory_156; // @[CPU.scala 52:20]
  reg [31:0] DMemory_157; // @[CPU.scala 52:20]
  reg [31:0] DMemory_158; // @[CPU.scala 52:20]
  reg [31:0] DMemory_159; // @[CPU.scala 52:20]
  reg [31:0] DMemory_160; // @[CPU.scala 52:20]
  reg [31:0] DMemory_161; // @[CPU.scala 52:20]
  reg [31:0] DMemory_162; // @[CPU.scala 52:20]
  reg [31:0] DMemory_163; // @[CPU.scala 52:20]
  reg [31:0] DMemory_164; // @[CPU.scala 52:20]
  reg [31:0] DMemory_165; // @[CPU.scala 52:20]
  reg [31:0] DMemory_166; // @[CPU.scala 52:20]
  reg [31:0] DMemory_167; // @[CPU.scala 52:20]
  reg [31:0] DMemory_168; // @[CPU.scala 52:20]
  reg [31:0] DMemory_169; // @[CPU.scala 52:20]
  reg [31:0] DMemory_170; // @[CPU.scala 52:20]
  reg [31:0] DMemory_171; // @[CPU.scala 52:20]
  reg [31:0] DMemory_172; // @[CPU.scala 52:20]
  reg [31:0] DMemory_173; // @[CPU.scala 52:20]
  reg [31:0] DMemory_174; // @[CPU.scala 52:20]
  reg [31:0] DMemory_175; // @[CPU.scala 52:20]
  reg [31:0] DMemory_176; // @[CPU.scala 52:20]
  reg [31:0] DMemory_177; // @[CPU.scala 52:20]
  reg [31:0] DMemory_178; // @[CPU.scala 52:20]
  reg [31:0] DMemory_179; // @[CPU.scala 52:20]
  reg [31:0] DMemory_180; // @[CPU.scala 52:20]
  reg [31:0] DMemory_181; // @[CPU.scala 52:20]
  reg [31:0] DMemory_182; // @[CPU.scala 52:20]
  reg [31:0] DMemory_183; // @[CPU.scala 52:20]
  reg [31:0] DMemory_184; // @[CPU.scala 52:20]
  reg [31:0] DMemory_185; // @[CPU.scala 52:20]
  reg [31:0] DMemory_186; // @[CPU.scala 52:20]
  reg [31:0] DMemory_187; // @[CPU.scala 52:20]
  reg [31:0] DMemory_188; // @[CPU.scala 52:20]
  reg [31:0] DMemory_189; // @[CPU.scala 52:20]
  reg [31:0] DMemory_190; // @[CPU.scala 52:20]
  reg [31:0] DMemory_191; // @[CPU.scala 52:20]
  reg [31:0] DMemory_192; // @[CPU.scala 52:20]
  reg [31:0] DMemory_193; // @[CPU.scala 52:20]
  reg [31:0] DMemory_194; // @[CPU.scala 52:20]
  reg [31:0] DMemory_195; // @[CPU.scala 52:20]
  reg [31:0] DMemory_196; // @[CPU.scala 52:20]
  reg [31:0] DMemory_197; // @[CPU.scala 52:20]
  reg [31:0] DMemory_198; // @[CPU.scala 52:20]
  reg [31:0] DMemory_199; // @[CPU.scala 52:20]
  reg [31:0] DMemory_200; // @[CPU.scala 52:20]
  reg [31:0] DMemory_201; // @[CPU.scala 52:20]
  reg [31:0] DMemory_202; // @[CPU.scala 52:20]
  reg [31:0] DMemory_203; // @[CPU.scala 52:20]
  reg [31:0] DMemory_204; // @[CPU.scala 52:20]
  reg [31:0] DMemory_205; // @[CPU.scala 52:20]
  reg [31:0] DMemory_206; // @[CPU.scala 52:20]
  reg [31:0] DMemory_207; // @[CPU.scala 52:20]
  reg [31:0] DMemory_208; // @[CPU.scala 52:20]
  reg [31:0] DMemory_209; // @[CPU.scala 52:20]
  reg [31:0] DMemory_210; // @[CPU.scala 52:20]
  reg [31:0] DMemory_211; // @[CPU.scala 52:20]
  reg [31:0] DMemory_212; // @[CPU.scala 52:20]
  reg [31:0] DMemory_213; // @[CPU.scala 52:20]
  reg [31:0] DMemory_214; // @[CPU.scala 52:20]
  reg [31:0] DMemory_215; // @[CPU.scala 52:20]
  reg [31:0] DMemory_216; // @[CPU.scala 52:20]
  reg [31:0] DMemory_217; // @[CPU.scala 52:20]
  reg [31:0] DMemory_218; // @[CPU.scala 52:20]
  reg [31:0] DMemory_219; // @[CPU.scala 52:20]
  reg [31:0] DMemory_220; // @[CPU.scala 52:20]
  reg [31:0] DMemory_221; // @[CPU.scala 52:20]
  reg [31:0] DMemory_222; // @[CPU.scala 52:20]
  reg [31:0] DMemory_223; // @[CPU.scala 52:20]
  reg [31:0] DMemory_224; // @[CPU.scala 52:20]
  reg [31:0] DMemory_225; // @[CPU.scala 52:20]
  reg [31:0] DMemory_226; // @[CPU.scala 52:20]
  reg [31:0] DMemory_227; // @[CPU.scala 52:20]
  reg [31:0] DMemory_228; // @[CPU.scala 52:20]
  reg [31:0] DMemory_229; // @[CPU.scala 52:20]
  reg [31:0] DMemory_230; // @[CPU.scala 52:20]
  reg [31:0] DMemory_231; // @[CPU.scala 52:20]
  reg [31:0] DMemory_232; // @[CPU.scala 52:20]
  reg [31:0] DMemory_233; // @[CPU.scala 52:20]
  reg [31:0] DMemory_234; // @[CPU.scala 52:20]
  reg [31:0] DMemory_235; // @[CPU.scala 52:20]
  reg [31:0] DMemory_236; // @[CPU.scala 52:20]
  reg [31:0] DMemory_237; // @[CPU.scala 52:20]
  reg [31:0] DMemory_238; // @[CPU.scala 52:20]
  reg [31:0] DMemory_239; // @[CPU.scala 52:20]
  reg [31:0] DMemory_240; // @[CPU.scala 52:20]
  reg [31:0] DMemory_241; // @[CPU.scala 52:20]
  reg [31:0] DMemory_242; // @[CPU.scala 52:20]
  reg [31:0] DMemory_243; // @[CPU.scala 52:20]
  reg [31:0] DMemory_244; // @[CPU.scala 52:20]
  reg [31:0] DMemory_245; // @[CPU.scala 52:20]
  reg [31:0] DMemory_246; // @[CPU.scala 52:20]
  reg [31:0] DMemory_247; // @[CPU.scala 52:20]
  reg [31:0] DMemory_248; // @[CPU.scala 52:20]
  reg [31:0] DMemory_249; // @[CPU.scala 52:20]
  reg [31:0] DMemory_250; // @[CPU.scala 52:20]
  reg [31:0] DMemory_251; // @[CPU.scala 52:20]
  reg [31:0] DMemory_252; // @[CPU.scala 52:20]
  reg [31:0] DMemory_253; // @[CPU.scala 52:20]
  reg [31:0] DMemory_254; // @[CPU.scala 52:20]
  reg [31:0] DMemory_255; // @[CPU.scala 52:20]
  reg [31:0] DMemory_256; // @[CPU.scala 52:20]
  reg [31:0] DMemory_257; // @[CPU.scala 52:20]
  reg [31:0] DMemory_258; // @[CPU.scala 52:20]
  reg [31:0] DMemory_259; // @[CPU.scala 52:20]
  reg [31:0] DMemory_260; // @[CPU.scala 52:20]
  reg [31:0] DMemory_261; // @[CPU.scala 52:20]
  reg [31:0] DMemory_262; // @[CPU.scala 52:20]
  reg [31:0] DMemory_263; // @[CPU.scala 52:20]
  reg [31:0] DMemory_264; // @[CPU.scala 52:20]
  reg [31:0] DMemory_265; // @[CPU.scala 52:20]
  reg [31:0] DMemory_266; // @[CPU.scala 52:20]
  reg [31:0] DMemory_267; // @[CPU.scala 52:20]
  reg [31:0] DMemory_268; // @[CPU.scala 52:20]
  reg [31:0] DMemory_269; // @[CPU.scala 52:20]
  reg [31:0] DMemory_270; // @[CPU.scala 52:20]
  reg [31:0] DMemory_271; // @[CPU.scala 52:20]
  reg [31:0] DMemory_272; // @[CPU.scala 52:20]
  reg [31:0] DMemory_273; // @[CPU.scala 52:20]
  reg [31:0] DMemory_274; // @[CPU.scala 52:20]
  reg [31:0] DMemory_275; // @[CPU.scala 52:20]
  reg [31:0] DMemory_276; // @[CPU.scala 52:20]
  reg [31:0] DMemory_277; // @[CPU.scala 52:20]
  reg [31:0] DMemory_278; // @[CPU.scala 52:20]
  reg [31:0] DMemory_279; // @[CPU.scala 52:20]
  reg [31:0] DMemory_280; // @[CPU.scala 52:20]
  reg [31:0] DMemory_281; // @[CPU.scala 52:20]
  reg [31:0] DMemory_282; // @[CPU.scala 52:20]
  reg [31:0] DMemory_283; // @[CPU.scala 52:20]
  reg [31:0] DMemory_284; // @[CPU.scala 52:20]
  reg [31:0] DMemory_285; // @[CPU.scala 52:20]
  reg [31:0] DMemory_286; // @[CPU.scala 52:20]
  reg [31:0] DMemory_287; // @[CPU.scala 52:20]
  reg [31:0] DMemory_288; // @[CPU.scala 52:20]
  reg [31:0] DMemory_289; // @[CPU.scala 52:20]
  reg [31:0] DMemory_290; // @[CPU.scala 52:20]
  reg [31:0] DMemory_291; // @[CPU.scala 52:20]
  reg [31:0] DMemory_292; // @[CPU.scala 52:20]
  reg [31:0] DMemory_293; // @[CPU.scala 52:20]
  reg [31:0] DMemory_294; // @[CPU.scala 52:20]
  reg [31:0] DMemory_295; // @[CPU.scala 52:20]
  reg [31:0] DMemory_296; // @[CPU.scala 52:20]
  reg [31:0] DMemory_297; // @[CPU.scala 52:20]
  reg [31:0] DMemory_298; // @[CPU.scala 52:20]
  reg [31:0] DMemory_299; // @[CPU.scala 52:20]
  reg [31:0] DMemory_300; // @[CPU.scala 52:20]
  reg [31:0] DMemory_301; // @[CPU.scala 52:20]
  reg [31:0] DMemory_302; // @[CPU.scala 52:20]
  reg [31:0] DMemory_303; // @[CPU.scala 52:20]
  reg [31:0] DMemory_304; // @[CPU.scala 52:20]
  reg [31:0] DMemory_305; // @[CPU.scala 52:20]
  reg [31:0] DMemory_306; // @[CPU.scala 52:20]
  reg [31:0] DMemory_307; // @[CPU.scala 52:20]
  reg [31:0] DMemory_308; // @[CPU.scala 52:20]
  reg [31:0] DMemory_309; // @[CPU.scala 52:20]
  reg [31:0] DMemory_310; // @[CPU.scala 52:20]
  reg [31:0] DMemory_311; // @[CPU.scala 52:20]
  reg [31:0] DMemory_312; // @[CPU.scala 52:20]
  reg [31:0] DMemory_313; // @[CPU.scala 52:20]
  reg [31:0] DMemory_314; // @[CPU.scala 52:20]
  reg [31:0] DMemory_315; // @[CPU.scala 52:20]
  reg [31:0] DMemory_316; // @[CPU.scala 52:20]
  reg [31:0] DMemory_317; // @[CPU.scala 52:20]
  reg [31:0] DMemory_318; // @[CPU.scala 52:20]
  reg [31:0] DMemory_319; // @[CPU.scala 52:20]
  reg [31:0] DMemory_320; // @[CPU.scala 52:20]
  reg [31:0] DMemory_321; // @[CPU.scala 52:20]
  reg [31:0] DMemory_322; // @[CPU.scala 52:20]
  reg [31:0] DMemory_323; // @[CPU.scala 52:20]
  reg [31:0] DMemory_324; // @[CPU.scala 52:20]
  reg [31:0] DMemory_325; // @[CPU.scala 52:20]
  reg [31:0] DMemory_326; // @[CPU.scala 52:20]
  reg [31:0] DMemory_327; // @[CPU.scala 52:20]
  reg [31:0] DMemory_328; // @[CPU.scala 52:20]
  reg [31:0] DMemory_329; // @[CPU.scala 52:20]
  reg [31:0] DMemory_330; // @[CPU.scala 52:20]
  reg [31:0] DMemory_331; // @[CPU.scala 52:20]
  reg [31:0] DMemory_332; // @[CPU.scala 52:20]
  reg [31:0] DMemory_333; // @[CPU.scala 52:20]
  reg [31:0] DMemory_334; // @[CPU.scala 52:20]
  reg [31:0] DMemory_335; // @[CPU.scala 52:20]
  reg [31:0] DMemory_336; // @[CPU.scala 52:20]
  reg [31:0] DMemory_337; // @[CPU.scala 52:20]
  reg [31:0] DMemory_338; // @[CPU.scala 52:20]
  reg [31:0] DMemory_339; // @[CPU.scala 52:20]
  reg [31:0] DMemory_340; // @[CPU.scala 52:20]
  reg [31:0] DMemory_341; // @[CPU.scala 52:20]
  reg [31:0] DMemory_342; // @[CPU.scala 52:20]
  reg [31:0] DMemory_343; // @[CPU.scala 52:20]
  reg [31:0] DMemory_344; // @[CPU.scala 52:20]
  reg [31:0] DMemory_345; // @[CPU.scala 52:20]
  reg [31:0] DMemory_346; // @[CPU.scala 52:20]
  reg [31:0] DMemory_347; // @[CPU.scala 52:20]
  reg [31:0] DMemory_348; // @[CPU.scala 52:20]
  reg [31:0] DMemory_349; // @[CPU.scala 52:20]
  reg [31:0] DMemory_350; // @[CPU.scala 52:20]
  reg [31:0] DMemory_351; // @[CPU.scala 52:20]
  reg [31:0] DMemory_352; // @[CPU.scala 52:20]
  reg [31:0] DMemory_353; // @[CPU.scala 52:20]
  reg [31:0] DMemory_354; // @[CPU.scala 52:20]
  reg [31:0] DMemory_355; // @[CPU.scala 52:20]
  reg [31:0] DMemory_356; // @[CPU.scala 52:20]
  reg [31:0] DMemory_357; // @[CPU.scala 52:20]
  reg [31:0] DMemory_358; // @[CPU.scala 52:20]
  reg [31:0] DMemory_359; // @[CPU.scala 52:20]
  reg [31:0] DMemory_360; // @[CPU.scala 52:20]
  reg [31:0] DMemory_361; // @[CPU.scala 52:20]
  reg [31:0] DMemory_362; // @[CPU.scala 52:20]
  reg [31:0] DMemory_363; // @[CPU.scala 52:20]
  reg [31:0] DMemory_364; // @[CPU.scala 52:20]
  reg [31:0] DMemory_365; // @[CPU.scala 52:20]
  reg [31:0] DMemory_366; // @[CPU.scala 52:20]
  reg [31:0] DMemory_367; // @[CPU.scala 52:20]
  reg [31:0] DMemory_368; // @[CPU.scala 52:20]
  reg [31:0] DMemory_369; // @[CPU.scala 52:20]
  reg [31:0] DMemory_370; // @[CPU.scala 52:20]
  reg [31:0] DMemory_371; // @[CPU.scala 52:20]
  reg [31:0] DMemory_372; // @[CPU.scala 52:20]
  reg [31:0] DMemory_373; // @[CPU.scala 52:20]
  reg [31:0] DMemory_374; // @[CPU.scala 52:20]
  reg [31:0] DMemory_375; // @[CPU.scala 52:20]
  reg [31:0] DMemory_376; // @[CPU.scala 52:20]
  reg [31:0] DMemory_377; // @[CPU.scala 52:20]
  reg [31:0] DMemory_378; // @[CPU.scala 52:20]
  reg [31:0] DMemory_379; // @[CPU.scala 52:20]
  reg [31:0] DMemory_380; // @[CPU.scala 52:20]
  reg [31:0] DMemory_381; // @[CPU.scala 52:20]
  reg [31:0] DMemory_382; // @[CPU.scala 52:20]
  reg [31:0] DMemory_383; // @[CPU.scala 52:20]
  reg [31:0] DMemory_384; // @[CPU.scala 52:20]
  reg [31:0] DMemory_385; // @[CPU.scala 52:20]
  reg [31:0] DMemory_386; // @[CPU.scala 52:20]
  reg [31:0] DMemory_387; // @[CPU.scala 52:20]
  reg [31:0] DMemory_388; // @[CPU.scala 52:20]
  reg [31:0] DMemory_389; // @[CPU.scala 52:20]
  reg [31:0] DMemory_390; // @[CPU.scala 52:20]
  reg [31:0] DMemory_391; // @[CPU.scala 52:20]
  reg [31:0] DMemory_392; // @[CPU.scala 52:20]
  reg [31:0] DMemory_393; // @[CPU.scala 52:20]
  reg [31:0] DMemory_394; // @[CPU.scala 52:20]
  reg [31:0] DMemory_395; // @[CPU.scala 52:20]
  reg [31:0] DMemory_396; // @[CPU.scala 52:20]
  reg [31:0] DMemory_397; // @[CPU.scala 52:20]
  reg [31:0] DMemory_398; // @[CPU.scala 52:20]
  reg [31:0] DMemory_399; // @[CPU.scala 52:20]
  reg [31:0] DMemory_400; // @[CPU.scala 52:20]
  reg [31:0] DMemory_401; // @[CPU.scala 52:20]
  reg [31:0] DMemory_402; // @[CPU.scala 52:20]
  reg [31:0] DMemory_403; // @[CPU.scala 52:20]
  reg [31:0] DMemory_404; // @[CPU.scala 52:20]
  reg [31:0] DMemory_405; // @[CPU.scala 52:20]
  reg [31:0] DMemory_406; // @[CPU.scala 52:20]
  reg [31:0] DMemory_407; // @[CPU.scala 52:20]
  reg [31:0] DMemory_408; // @[CPU.scala 52:20]
  reg [31:0] DMemory_409; // @[CPU.scala 52:20]
  reg [31:0] DMemory_410; // @[CPU.scala 52:20]
  reg [31:0] DMemory_411; // @[CPU.scala 52:20]
  reg [31:0] DMemory_412; // @[CPU.scala 52:20]
  reg [31:0] DMemory_413; // @[CPU.scala 52:20]
  reg [31:0] DMemory_414; // @[CPU.scala 52:20]
  reg [31:0] DMemory_415; // @[CPU.scala 52:20]
  reg [31:0] DMemory_416; // @[CPU.scala 52:20]
  reg [31:0] DMemory_417; // @[CPU.scala 52:20]
  reg [31:0] DMemory_418; // @[CPU.scala 52:20]
  reg [31:0] DMemory_419; // @[CPU.scala 52:20]
  reg [31:0] DMemory_420; // @[CPU.scala 52:20]
  reg [31:0] DMemory_421; // @[CPU.scala 52:20]
  reg [31:0] DMemory_422; // @[CPU.scala 52:20]
  reg [31:0] DMemory_423; // @[CPU.scala 52:20]
  reg [31:0] DMemory_424; // @[CPU.scala 52:20]
  reg [31:0] DMemory_425; // @[CPU.scala 52:20]
  reg [31:0] DMemory_426; // @[CPU.scala 52:20]
  reg [31:0] DMemory_427; // @[CPU.scala 52:20]
  reg [31:0] DMemory_428; // @[CPU.scala 52:20]
  reg [31:0] DMemory_429; // @[CPU.scala 52:20]
  reg [31:0] DMemory_430; // @[CPU.scala 52:20]
  reg [31:0] DMemory_431; // @[CPU.scala 52:20]
  reg [31:0] DMemory_432; // @[CPU.scala 52:20]
  reg [31:0] DMemory_433; // @[CPU.scala 52:20]
  reg [31:0] DMemory_434; // @[CPU.scala 52:20]
  reg [31:0] DMemory_435; // @[CPU.scala 52:20]
  reg [31:0] DMemory_436; // @[CPU.scala 52:20]
  reg [31:0] DMemory_437; // @[CPU.scala 52:20]
  reg [31:0] DMemory_438; // @[CPU.scala 52:20]
  reg [31:0] DMemory_439; // @[CPU.scala 52:20]
  reg [31:0] DMemory_440; // @[CPU.scala 52:20]
  reg [31:0] DMemory_441; // @[CPU.scala 52:20]
  reg [31:0] DMemory_442; // @[CPU.scala 52:20]
  reg [31:0] DMemory_443; // @[CPU.scala 52:20]
  reg [31:0] DMemory_444; // @[CPU.scala 52:20]
  reg [31:0] DMemory_445; // @[CPU.scala 52:20]
  reg [31:0] DMemory_446; // @[CPU.scala 52:20]
  reg [31:0] DMemory_447; // @[CPU.scala 52:20]
  reg [31:0] DMemory_448; // @[CPU.scala 52:20]
  reg [31:0] DMemory_449; // @[CPU.scala 52:20]
  reg [31:0] DMemory_450; // @[CPU.scala 52:20]
  reg [31:0] DMemory_451; // @[CPU.scala 52:20]
  reg [31:0] DMemory_452; // @[CPU.scala 52:20]
  reg [31:0] DMemory_453; // @[CPU.scala 52:20]
  reg [31:0] DMemory_454; // @[CPU.scala 52:20]
  reg [31:0] DMemory_455; // @[CPU.scala 52:20]
  reg [31:0] DMemory_456; // @[CPU.scala 52:20]
  reg [31:0] DMemory_457; // @[CPU.scala 52:20]
  reg [31:0] DMemory_458; // @[CPU.scala 52:20]
  reg [31:0] DMemory_459; // @[CPU.scala 52:20]
  reg [31:0] DMemory_460; // @[CPU.scala 52:20]
  reg [31:0] DMemory_461; // @[CPU.scala 52:20]
  reg [31:0] DMemory_462; // @[CPU.scala 52:20]
  reg [31:0] DMemory_463; // @[CPU.scala 52:20]
  reg [31:0] DMemory_464; // @[CPU.scala 52:20]
  reg [31:0] DMemory_465; // @[CPU.scala 52:20]
  reg [31:0] DMemory_466; // @[CPU.scala 52:20]
  reg [31:0] DMemory_467; // @[CPU.scala 52:20]
  reg [31:0] DMemory_468; // @[CPU.scala 52:20]
  reg [31:0] DMemory_469; // @[CPU.scala 52:20]
  reg [31:0] DMemory_470; // @[CPU.scala 52:20]
  reg [31:0] DMemory_471; // @[CPU.scala 52:20]
  reg [31:0] DMemory_472; // @[CPU.scala 52:20]
  reg [31:0] DMemory_473; // @[CPU.scala 52:20]
  reg [31:0] DMemory_474; // @[CPU.scala 52:20]
  reg [31:0] DMemory_475; // @[CPU.scala 52:20]
  reg [31:0] DMemory_476; // @[CPU.scala 52:20]
  reg [31:0] DMemory_477; // @[CPU.scala 52:20]
  reg [31:0] DMemory_478; // @[CPU.scala 52:20]
  reg [31:0] DMemory_479; // @[CPU.scala 52:20]
  reg [31:0] DMemory_480; // @[CPU.scala 52:20]
  reg [31:0] DMemory_481; // @[CPU.scala 52:20]
  reg [31:0] DMemory_482; // @[CPU.scala 52:20]
  reg [31:0] DMemory_483; // @[CPU.scala 52:20]
  reg [31:0] DMemory_484; // @[CPU.scala 52:20]
  reg [31:0] DMemory_485; // @[CPU.scala 52:20]
  reg [31:0] DMemory_486; // @[CPU.scala 52:20]
  reg [31:0] DMemory_487; // @[CPU.scala 52:20]
  reg [31:0] DMemory_488; // @[CPU.scala 52:20]
  reg [31:0] DMemory_489; // @[CPU.scala 52:20]
  reg [31:0] DMemory_490; // @[CPU.scala 52:20]
  reg [31:0] DMemory_491; // @[CPU.scala 52:20]
  reg [31:0] DMemory_492; // @[CPU.scala 52:20]
  reg [31:0] DMemory_493; // @[CPU.scala 52:20]
  reg [31:0] DMemory_494; // @[CPU.scala 52:20]
  reg [31:0] DMemory_495; // @[CPU.scala 52:20]
  reg [31:0] DMemory_496; // @[CPU.scala 52:20]
  reg [31:0] DMemory_497; // @[CPU.scala 52:20]
  reg [31:0] DMemory_498; // @[CPU.scala 52:20]
  reg [31:0] DMemory_499; // @[CPU.scala 52:20]
  reg [31:0] DMemory_500; // @[CPU.scala 52:20]
  reg [31:0] DMemory_501; // @[CPU.scala 52:20]
  reg [31:0] DMemory_502; // @[CPU.scala 52:20]
  reg [31:0] DMemory_503; // @[CPU.scala 52:20]
  reg [31:0] DMemory_504; // @[CPU.scala 52:20]
  reg [31:0] DMemory_505; // @[CPU.scala 52:20]
  reg [31:0] DMemory_506; // @[CPU.scala 52:20]
  reg [31:0] DMemory_507; // @[CPU.scala 52:20]
  reg [31:0] DMemory_508; // @[CPU.scala 52:20]
  reg [31:0] DMemory_509; // @[CPU.scala 52:20]
  reg [31:0] DMemory_510; // @[CPU.scala 52:20]
  reg [31:0] DMemory_511; // @[CPU.scala 52:20]
  reg [31:0] DMemory_512; // @[CPU.scala 52:20]
  reg [31:0] DMemory_513; // @[CPU.scala 52:20]
  reg [31:0] DMemory_514; // @[CPU.scala 52:20]
  reg [31:0] DMemory_515; // @[CPU.scala 52:20]
  reg [31:0] DMemory_516; // @[CPU.scala 52:20]
  reg [31:0] DMemory_517; // @[CPU.scala 52:20]
  reg [31:0] DMemory_518; // @[CPU.scala 52:20]
  reg [31:0] DMemory_519; // @[CPU.scala 52:20]
  reg [31:0] DMemory_520; // @[CPU.scala 52:20]
  reg [31:0] DMemory_521; // @[CPU.scala 52:20]
  reg [31:0] DMemory_522; // @[CPU.scala 52:20]
  reg [31:0] DMemory_523; // @[CPU.scala 52:20]
  reg [31:0] DMemory_524; // @[CPU.scala 52:20]
  reg [31:0] DMemory_525; // @[CPU.scala 52:20]
  reg [31:0] DMemory_526; // @[CPU.scala 52:20]
  reg [31:0] DMemory_527; // @[CPU.scala 52:20]
  reg [31:0] DMemory_528; // @[CPU.scala 52:20]
  reg [31:0] DMemory_529; // @[CPU.scala 52:20]
  reg [31:0] DMemory_530; // @[CPU.scala 52:20]
  reg [31:0] DMemory_531; // @[CPU.scala 52:20]
  reg [31:0] DMemory_532; // @[CPU.scala 52:20]
  reg [31:0] DMemory_533; // @[CPU.scala 52:20]
  reg [31:0] DMemory_534; // @[CPU.scala 52:20]
  reg [31:0] DMemory_535; // @[CPU.scala 52:20]
  reg [31:0] DMemory_536; // @[CPU.scala 52:20]
  reg [31:0] DMemory_537; // @[CPU.scala 52:20]
  reg [31:0] DMemory_538; // @[CPU.scala 52:20]
  reg [31:0] DMemory_539; // @[CPU.scala 52:20]
  reg [31:0] DMemory_540; // @[CPU.scala 52:20]
  reg [31:0] DMemory_541; // @[CPU.scala 52:20]
  reg [31:0] DMemory_542; // @[CPU.scala 52:20]
  reg [31:0] DMemory_543; // @[CPU.scala 52:20]
  reg [31:0] DMemory_544; // @[CPU.scala 52:20]
  reg [31:0] DMemory_545; // @[CPU.scala 52:20]
  reg [31:0] DMemory_546; // @[CPU.scala 52:20]
  reg [31:0] DMemory_547; // @[CPU.scala 52:20]
  reg [31:0] DMemory_548; // @[CPU.scala 52:20]
  reg [31:0] DMemory_549; // @[CPU.scala 52:20]
  reg [31:0] DMemory_550; // @[CPU.scala 52:20]
  reg [31:0] DMemory_551; // @[CPU.scala 52:20]
  reg [31:0] DMemory_552; // @[CPU.scala 52:20]
  reg [31:0] DMemory_553; // @[CPU.scala 52:20]
  reg [31:0] DMemory_554; // @[CPU.scala 52:20]
  reg [31:0] DMemory_555; // @[CPU.scala 52:20]
  reg [31:0] DMemory_556; // @[CPU.scala 52:20]
  reg [31:0] DMemory_557; // @[CPU.scala 52:20]
  reg [31:0] DMemory_558; // @[CPU.scala 52:20]
  reg [31:0] DMemory_559; // @[CPU.scala 52:20]
  reg [31:0] DMemory_560; // @[CPU.scala 52:20]
  reg [31:0] DMemory_561; // @[CPU.scala 52:20]
  reg [31:0] DMemory_562; // @[CPU.scala 52:20]
  reg [31:0] DMemory_563; // @[CPU.scala 52:20]
  reg [31:0] DMemory_564; // @[CPU.scala 52:20]
  reg [31:0] DMemory_565; // @[CPU.scala 52:20]
  reg [31:0] DMemory_566; // @[CPU.scala 52:20]
  reg [31:0] DMemory_567; // @[CPU.scala 52:20]
  reg [31:0] DMemory_568; // @[CPU.scala 52:20]
  reg [31:0] DMemory_569; // @[CPU.scala 52:20]
  reg [31:0] DMemory_570; // @[CPU.scala 52:20]
  reg [31:0] DMemory_571; // @[CPU.scala 52:20]
  reg [31:0] DMemory_572; // @[CPU.scala 52:20]
  reg [31:0] DMemory_573; // @[CPU.scala 52:20]
  reg [31:0] DMemory_574; // @[CPU.scala 52:20]
  reg [31:0] DMemory_575; // @[CPU.scala 52:20]
  reg [31:0] DMemory_576; // @[CPU.scala 52:20]
  reg [31:0] DMemory_577; // @[CPU.scala 52:20]
  reg [31:0] DMemory_578; // @[CPU.scala 52:20]
  reg [31:0] DMemory_579; // @[CPU.scala 52:20]
  reg [31:0] DMemory_580; // @[CPU.scala 52:20]
  reg [31:0] DMemory_581; // @[CPU.scala 52:20]
  reg [31:0] DMemory_582; // @[CPU.scala 52:20]
  reg [31:0] DMemory_583; // @[CPU.scala 52:20]
  reg [31:0] DMemory_584; // @[CPU.scala 52:20]
  reg [31:0] DMemory_585; // @[CPU.scala 52:20]
  reg [31:0] DMemory_586; // @[CPU.scala 52:20]
  reg [31:0] DMemory_587; // @[CPU.scala 52:20]
  reg [31:0] DMemory_588; // @[CPU.scala 52:20]
  reg [31:0] DMemory_589; // @[CPU.scala 52:20]
  reg [31:0] DMemory_590; // @[CPU.scala 52:20]
  reg [31:0] DMemory_591; // @[CPU.scala 52:20]
  reg [31:0] DMemory_592; // @[CPU.scala 52:20]
  reg [31:0] DMemory_593; // @[CPU.scala 52:20]
  reg [31:0] DMemory_594; // @[CPU.scala 52:20]
  reg [31:0] DMemory_595; // @[CPU.scala 52:20]
  reg [31:0] DMemory_596; // @[CPU.scala 52:20]
  reg [31:0] DMemory_597; // @[CPU.scala 52:20]
  reg [31:0] DMemory_598; // @[CPU.scala 52:20]
  reg [31:0] DMemory_599; // @[CPU.scala 52:20]
  reg [31:0] DMemory_600; // @[CPU.scala 52:20]
  reg [31:0] DMemory_601; // @[CPU.scala 52:20]
  reg [31:0] DMemory_602; // @[CPU.scala 52:20]
  reg [31:0] DMemory_603; // @[CPU.scala 52:20]
  reg [31:0] DMemory_604; // @[CPU.scala 52:20]
  reg [31:0] DMemory_605; // @[CPU.scala 52:20]
  reg [31:0] DMemory_606; // @[CPU.scala 52:20]
  reg [31:0] DMemory_607; // @[CPU.scala 52:20]
  reg [31:0] DMemory_608; // @[CPU.scala 52:20]
  reg [31:0] DMemory_609; // @[CPU.scala 52:20]
  reg [31:0] DMemory_610; // @[CPU.scala 52:20]
  reg [31:0] DMemory_611; // @[CPU.scala 52:20]
  reg [31:0] DMemory_612; // @[CPU.scala 52:20]
  reg [31:0] DMemory_613; // @[CPU.scala 52:20]
  reg [31:0] DMemory_614; // @[CPU.scala 52:20]
  reg [31:0] DMemory_615; // @[CPU.scala 52:20]
  reg [31:0] DMemory_616; // @[CPU.scala 52:20]
  reg [31:0] DMemory_617; // @[CPU.scala 52:20]
  reg [31:0] DMemory_618; // @[CPU.scala 52:20]
  reg [31:0] DMemory_619; // @[CPU.scala 52:20]
  reg [31:0] DMemory_620; // @[CPU.scala 52:20]
  reg [31:0] DMemory_621; // @[CPU.scala 52:20]
  reg [31:0] DMemory_622; // @[CPU.scala 52:20]
  reg [31:0] DMemory_623; // @[CPU.scala 52:20]
  reg [31:0] DMemory_624; // @[CPU.scala 52:20]
  reg [31:0] DMemory_625; // @[CPU.scala 52:20]
  reg [31:0] DMemory_626; // @[CPU.scala 52:20]
  reg [31:0] DMemory_627; // @[CPU.scala 52:20]
  reg [31:0] DMemory_628; // @[CPU.scala 52:20]
  reg [31:0] DMemory_629; // @[CPU.scala 52:20]
  reg [31:0] DMemory_630; // @[CPU.scala 52:20]
  reg [31:0] DMemory_631; // @[CPU.scala 52:20]
  reg [31:0] DMemory_632; // @[CPU.scala 52:20]
  reg [31:0] DMemory_633; // @[CPU.scala 52:20]
  reg [31:0] DMemory_634; // @[CPU.scala 52:20]
  reg [31:0] DMemory_635; // @[CPU.scala 52:20]
  reg [31:0] DMemory_636; // @[CPU.scala 52:20]
  reg [31:0] DMemory_637; // @[CPU.scala 52:20]
  reg [31:0] DMemory_638; // @[CPU.scala 52:20]
  reg [31:0] DMemory_639; // @[CPU.scala 52:20]
  reg [31:0] DMemory_640; // @[CPU.scala 52:20]
  reg [31:0] DMemory_641; // @[CPU.scala 52:20]
  reg [31:0] DMemory_642; // @[CPU.scala 52:20]
  reg [31:0] DMemory_643; // @[CPU.scala 52:20]
  reg [31:0] DMemory_644; // @[CPU.scala 52:20]
  reg [31:0] DMemory_645; // @[CPU.scala 52:20]
  reg [31:0] DMemory_646; // @[CPU.scala 52:20]
  reg [31:0] DMemory_647; // @[CPU.scala 52:20]
  reg [31:0] DMemory_648; // @[CPU.scala 52:20]
  reg [31:0] DMemory_649; // @[CPU.scala 52:20]
  reg [31:0] DMemory_650; // @[CPU.scala 52:20]
  reg [31:0] DMemory_651; // @[CPU.scala 52:20]
  reg [31:0] DMemory_652; // @[CPU.scala 52:20]
  reg [31:0] DMemory_653; // @[CPU.scala 52:20]
  reg [31:0] DMemory_654; // @[CPU.scala 52:20]
  reg [31:0] DMemory_655; // @[CPU.scala 52:20]
  reg [31:0] DMemory_656; // @[CPU.scala 52:20]
  reg [31:0] DMemory_657; // @[CPU.scala 52:20]
  reg [31:0] DMemory_658; // @[CPU.scala 52:20]
  reg [31:0] DMemory_659; // @[CPU.scala 52:20]
  reg [31:0] DMemory_660; // @[CPU.scala 52:20]
  reg [31:0] DMemory_661; // @[CPU.scala 52:20]
  reg [31:0] DMemory_662; // @[CPU.scala 52:20]
  reg [31:0] DMemory_663; // @[CPU.scala 52:20]
  reg [31:0] DMemory_664; // @[CPU.scala 52:20]
  reg [31:0] DMemory_665; // @[CPU.scala 52:20]
  reg [31:0] DMemory_666; // @[CPU.scala 52:20]
  reg [31:0] DMemory_667; // @[CPU.scala 52:20]
  reg [31:0] DMemory_668; // @[CPU.scala 52:20]
  reg [31:0] DMemory_669; // @[CPU.scala 52:20]
  reg [31:0] DMemory_670; // @[CPU.scala 52:20]
  reg [31:0] DMemory_671; // @[CPU.scala 52:20]
  reg [31:0] DMemory_672; // @[CPU.scala 52:20]
  reg [31:0] DMemory_673; // @[CPU.scala 52:20]
  reg [31:0] DMemory_674; // @[CPU.scala 52:20]
  reg [31:0] DMemory_675; // @[CPU.scala 52:20]
  reg [31:0] DMemory_676; // @[CPU.scala 52:20]
  reg [31:0] DMemory_677; // @[CPU.scala 52:20]
  reg [31:0] DMemory_678; // @[CPU.scala 52:20]
  reg [31:0] DMemory_679; // @[CPU.scala 52:20]
  reg [31:0] DMemory_680; // @[CPU.scala 52:20]
  reg [31:0] DMemory_681; // @[CPU.scala 52:20]
  reg [31:0] DMemory_682; // @[CPU.scala 52:20]
  reg [31:0] DMemory_683; // @[CPU.scala 52:20]
  reg [31:0] DMemory_684; // @[CPU.scala 52:20]
  reg [31:0] DMemory_685; // @[CPU.scala 52:20]
  reg [31:0] DMemory_686; // @[CPU.scala 52:20]
  reg [31:0] DMemory_687; // @[CPU.scala 52:20]
  reg [31:0] DMemory_688; // @[CPU.scala 52:20]
  reg [31:0] DMemory_689; // @[CPU.scala 52:20]
  reg [31:0] DMemory_690; // @[CPU.scala 52:20]
  reg [31:0] DMemory_691; // @[CPU.scala 52:20]
  reg [31:0] DMemory_692; // @[CPU.scala 52:20]
  reg [31:0] DMemory_693; // @[CPU.scala 52:20]
  reg [31:0] DMemory_694; // @[CPU.scala 52:20]
  reg [31:0] DMemory_695; // @[CPU.scala 52:20]
  reg [31:0] DMemory_696; // @[CPU.scala 52:20]
  reg [31:0] DMemory_697; // @[CPU.scala 52:20]
  reg [31:0] DMemory_698; // @[CPU.scala 52:20]
  reg [31:0] DMemory_699; // @[CPU.scala 52:20]
  reg [31:0] DMemory_700; // @[CPU.scala 52:20]
  reg [31:0] DMemory_701; // @[CPU.scala 52:20]
  reg [31:0] DMemory_702; // @[CPU.scala 52:20]
  reg [31:0] DMemory_703; // @[CPU.scala 52:20]
  reg [31:0] DMemory_704; // @[CPU.scala 52:20]
  reg [31:0] DMemory_705; // @[CPU.scala 52:20]
  reg [31:0] DMemory_706; // @[CPU.scala 52:20]
  reg [31:0] DMemory_707; // @[CPU.scala 52:20]
  reg [31:0] DMemory_708; // @[CPU.scala 52:20]
  reg [31:0] DMemory_709; // @[CPU.scala 52:20]
  reg [31:0] DMemory_710; // @[CPU.scala 52:20]
  reg [31:0] DMemory_711; // @[CPU.scala 52:20]
  reg [31:0] DMemory_712; // @[CPU.scala 52:20]
  reg [31:0] DMemory_713; // @[CPU.scala 52:20]
  reg [31:0] DMemory_714; // @[CPU.scala 52:20]
  reg [31:0] DMemory_715; // @[CPU.scala 52:20]
  reg [31:0] DMemory_716; // @[CPU.scala 52:20]
  reg [31:0] DMemory_717; // @[CPU.scala 52:20]
  reg [31:0] DMemory_718; // @[CPU.scala 52:20]
  reg [31:0] DMemory_719; // @[CPU.scala 52:20]
  reg [31:0] DMemory_720; // @[CPU.scala 52:20]
  reg [31:0] DMemory_721; // @[CPU.scala 52:20]
  reg [31:0] DMemory_722; // @[CPU.scala 52:20]
  reg [31:0] DMemory_723; // @[CPU.scala 52:20]
  reg [31:0] DMemory_724; // @[CPU.scala 52:20]
  reg [31:0] DMemory_725; // @[CPU.scala 52:20]
  reg [31:0] DMemory_726; // @[CPU.scala 52:20]
  reg [31:0] DMemory_727; // @[CPU.scala 52:20]
  reg [31:0] DMemory_728; // @[CPU.scala 52:20]
  reg [31:0] DMemory_729; // @[CPU.scala 52:20]
  reg [31:0] DMemory_730; // @[CPU.scala 52:20]
  reg [31:0] DMemory_731; // @[CPU.scala 52:20]
  reg [31:0] DMemory_732; // @[CPU.scala 52:20]
  reg [31:0] DMemory_733; // @[CPU.scala 52:20]
  reg [31:0] DMemory_734; // @[CPU.scala 52:20]
  reg [31:0] DMemory_735; // @[CPU.scala 52:20]
  reg [31:0] DMemory_736; // @[CPU.scala 52:20]
  reg [31:0] DMemory_737; // @[CPU.scala 52:20]
  reg [31:0] DMemory_738; // @[CPU.scala 52:20]
  reg [31:0] DMemory_739; // @[CPU.scala 52:20]
  reg [31:0] DMemory_740; // @[CPU.scala 52:20]
  reg [31:0] DMemory_741; // @[CPU.scala 52:20]
  reg [31:0] DMemory_742; // @[CPU.scala 52:20]
  reg [31:0] DMemory_743; // @[CPU.scala 52:20]
  reg [31:0] DMemory_744; // @[CPU.scala 52:20]
  reg [31:0] DMemory_745; // @[CPU.scala 52:20]
  reg [31:0] DMemory_746; // @[CPU.scala 52:20]
  reg [31:0] DMemory_747; // @[CPU.scala 52:20]
  reg [31:0] DMemory_748; // @[CPU.scala 52:20]
  reg [31:0] DMemory_749; // @[CPU.scala 52:20]
  reg [31:0] DMemory_750; // @[CPU.scala 52:20]
  reg [31:0] DMemory_751; // @[CPU.scala 52:20]
  reg [31:0] DMemory_752; // @[CPU.scala 52:20]
  reg [31:0] DMemory_753; // @[CPU.scala 52:20]
  reg [31:0] DMemory_754; // @[CPU.scala 52:20]
  reg [31:0] DMemory_755; // @[CPU.scala 52:20]
  reg [31:0] DMemory_756; // @[CPU.scala 52:20]
  reg [31:0] DMemory_757; // @[CPU.scala 52:20]
  reg [31:0] DMemory_758; // @[CPU.scala 52:20]
  reg [31:0] DMemory_759; // @[CPU.scala 52:20]
  reg [31:0] DMemory_760; // @[CPU.scala 52:20]
  reg [31:0] DMemory_761; // @[CPU.scala 52:20]
  reg [31:0] DMemory_762; // @[CPU.scala 52:20]
  reg [31:0] DMemory_763; // @[CPU.scala 52:20]
  reg [31:0] DMemory_764; // @[CPU.scala 52:20]
  reg [31:0] DMemory_765; // @[CPU.scala 52:20]
  reg [31:0] DMemory_766; // @[CPU.scala 52:20]
  reg [31:0] DMemory_767; // @[CPU.scala 52:20]
  reg [31:0] DMemory_768; // @[CPU.scala 52:20]
  reg [31:0] DMemory_769; // @[CPU.scala 52:20]
  reg [31:0] DMemory_770; // @[CPU.scala 52:20]
  reg [31:0] DMemory_771; // @[CPU.scala 52:20]
  reg [31:0] DMemory_772; // @[CPU.scala 52:20]
  reg [31:0] DMemory_773; // @[CPU.scala 52:20]
  reg [31:0] DMemory_774; // @[CPU.scala 52:20]
  reg [31:0] DMemory_775; // @[CPU.scala 52:20]
  reg [31:0] DMemory_776; // @[CPU.scala 52:20]
  reg [31:0] DMemory_777; // @[CPU.scala 52:20]
  reg [31:0] DMemory_778; // @[CPU.scala 52:20]
  reg [31:0] DMemory_779; // @[CPU.scala 52:20]
  reg [31:0] DMemory_780; // @[CPU.scala 52:20]
  reg [31:0] DMemory_781; // @[CPU.scala 52:20]
  reg [31:0] DMemory_782; // @[CPU.scala 52:20]
  reg [31:0] DMemory_783; // @[CPU.scala 52:20]
  reg [31:0] DMemory_784; // @[CPU.scala 52:20]
  reg [31:0] DMemory_785; // @[CPU.scala 52:20]
  reg [31:0] DMemory_786; // @[CPU.scala 52:20]
  reg [31:0] DMemory_787; // @[CPU.scala 52:20]
  reg [31:0] DMemory_788; // @[CPU.scala 52:20]
  reg [31:0] DMemory_789; // @[CPU.scala 52:20]
  reg [31:0] DMemory_790; // @[CPU.scala 52:20]
  reg [31:0] DMemory_791; // @[CPU.scala 52:20]
  reg [31:0] DMemory_792; // @[CPU.scala 52:20]
  reg [31:0] DMemory_793; // @[CPU.scala 52:20]
  reg [31:0] DMemory_794; // @[CPU.scala 52:20]
  reg [31:0] DMemory_795; // @[CPU.scala 52:20]
  reg [31:0] DMemory_796; // @[CPU.scala 52:20]
  reg [31:0] DMemory_797; // @[CPU.scala 52:20]
  reg [31:0] DMemory_798; // @[CPU.scala 52:20]
  reg [31:0] DMemory_799; // @[CPU.scala 52:20]
  reg [31:0] DMemory_800; // @[CPU.scala 52:20]
  reg [31:0] DMemory_801; // @[CPU.scala 52:20]
  reg [31:0] DMemory_802; // @[CPU.scala 52:20]
  reg [31:0] DMemory_803; // @[CPU.scala 52:20]
  reg [31:0] DMemory_804; // @[CPU.scala 52:20]
  reg [31:0] DMemory_805; // @[CPU.scala 52:20]
  reg [31:0] DMemory_806; // @[CPU.scala 52:20]
  reg [31:0] DMemory_807; // @[CPU.scala 52:20]
  reg [31:0] DMemory_808; // @[CPU.scala 52:20]
  reg [31:0] DMemory_809; // @[CPU.scala 52:20]
  reg [31:0] DMemory_810; // @[CPU.scala 52:20]
  reg [31:0] DMemory_811; // @[CPU.scala 52:20]
  reg [31:0] DMemory_812; // @[CPU.scala 52:20]
  reg [31:0] DMemory_813; // @[CPU.scala 52:20]
  reg [31:0] DMemory_814; // @[CPU.scala 52:20]
  reg [31:0] DMemory_815; // @[CPU.scala 52:20]
  reg [31:0] DMemory_816; // @[CPU.scala 52:20]
  reg [31:0] DMemory_817; // @[CPU.scala 52:20]
  reg [31:0] DMemory_818; // @[CPU.scala 52:20]
  reg [31:0] DMemory_819; // @[CPU.scala 52:20]
  reg [31:0] DMemory_820; // @[CPU.scala 52:20]
  reg [31:0] DMemory_821; // @[CPU.scala 52:20]
  reg [31:0] DMemory_822; // @[CPU.scala 52:20]
  reg [31:0] DMemory_823; // @[CPU.scala 52:20]
  reg [31:0] DMemory_824; // @[CPU.scala 52:20]
  reg [31:0] DMemory_825; // @[CPU.scala 52:20]
  reg [31:0] DMemory_826; // @[CPU.scala 52:20]
  reg [31:0] DMemory_827; // @[CPU.scala 52:20]
  reg [31:0] DMemory_828; // @[CPU.scala 52:20]
  reg [31:0] DMemory_829; // @[CPU.scala 52:20]
  reg [31:0] DMemory_830; // @[CPU.scala 52:20]
  reg [31:0] DMemory_831; // @[CPU.scala 52:20]
  reg [31:0] DMemory_832; // @[CPU.scala 52:20]
  reg [31:0] DMemory_833; // @[CPU.scala 52:20]
  reg [31:0] DMemory_834; // @[CPU.scala 52:20]
  reg [31:0] DMemory_835; // @[CPU.scala 52:20]
  reg [31:0] DMemory_836; // @[CPU.scala 52:20]
  reg [31:0] DMemory_837; // @[CPU.scala 52:20]
  reg [31:0] DMemory_838; // @[CPU.scala 52:20]
  reg [31:0] DMemory_839; // @[CPU.scala 52:20]
  reg [31:0] DMemory_840; // @[CPU.scala 52:20]
  reg [31:0] DMemory_841; // @[CPU.scala 52:20]
  reg [31:0] DMemory_842; // @[CPU.scala 52:20]
  reg [31:0] DMemory_843; // @[CPU.scala 52:20]
  reg [31:0] DMemory_844; // @[CPU.scala 52:20]
  reg [31:0] DMemory_845; // @[CPU.scala 52:20]
  reg [31:0] DMemory_846; // @[CPU.scala 52:20]
  reg [31:0] DMemory_847; // @[CPU.scala 52:20]
  reg [31:0] DMemory_848; // @[CPU.scala 52:20]
  reg [31:0] DMemory_849; // @[CPU.scala 52:20]
  reg [31:0] DMemory_850; // @[CPU.scala 52:20]
  reg [31:0] DMemory_851; // @[CPU.scala 52:20]
  reg [31:0] DMemory_852; // @[CPU.scala 52:20]
  reg [31:0] DMemory_853; // @[CPU.scala 52:20]
  reg [31:0] DMemory_854; // @[CPU.scala 52:20]
  reg [31:0] DMemory_855; // @[CPU.scala 52:20]
  reg [31:0] DMemory_856; // @[CPU.scala 52:20]
  reg [31:0] DMemory_857; // @[CPU.scala 52:20]
  reg [31:0] DMemory_858; // @[CPU.scala 52:20]
  reg [31:0] DMemory_859; // @[CPU.scala 52:20]
  reg [31:0] DMemory_860; // @[CPU.scala 52:20]
  reg [31:0] DMemory_861; // @[CPU.scala 52:20]
  reg [31:0] DMemory_862; // @[CPU.scala 52:20]
  reg [31:0] DMemory_863; // @[CPU.scala 52:20]
  reg [31:0] DMemory_864; // @[CPU.scala 52:20]
  reg [31:0] DMemory_865; // @[CPU.scala 52:20]
  reg [31:0] DMemory_866; // @[CPU.scala 52:20]
  reg [31:0] DMemory_867; // @[CPU.scala 52:20]
  reg [31:0] DMemory_868; // @[CPU.scala 52:20]
  reg [31:0] DMemory_869; // @[CPU.scala 52:20]
  reg [31:0] DMemory_870; // @[CPU.scala 52:20]
  reg [31:0] DMemory_871; // @[CPU.scala 52:20]
  reg [31:0] DMemory_872; // @[CPU.scala 52:20]
  reg [31:0] DMemory_873; // @[CPU.scala 52:20]
  reg [31:0] DMemory_874; // @[CPU.scala 52:20]
  reg [31:0] DMemory_875; // @[CPU.scala 52:20]
  reg [31:0] DMemory_876; // @[CPU.scala 52:20]
  reg [31:0] DMemory_877; // @[CPU.scala 52:20]
  reg [31:0] DMemory_878; // @[CPU.scala 52:20]
  reg [31:0] DMemory_879; // @[CPU.scala 52:20]
  reg [31:0] DMemory_880; // @[CPU.scala 52:20]
  reg [31:0] DMemory_881; // @[CPU.scala 52:20]
  reg [31:0] DMemory_882; // @[CPU.scala 52:20]
  reg [31:0] DMemory_883; // @[CPU.scala 52:20]
  reg [31:0] DMemory_884; // @[CPU.scala 52:20]
  reg [31:0] DMemory_885; // @[CPU.scala 52:20]
  reg [31:0] DMemory_886; // @[CPU.scala 52:20]
  reg [31:0] DMemory_887; // @[CPU.scala 52:20]
  reg [31:0] DMemory_888; // @[CPU.scala 52:20]
  reg [31:0] DMemory_889; // @[CPU.scala 52:20]
  reg [31:0] DMemory_890; // @[CPU.scala 52:20]
  reg [31:0] DMemory_891; // @[CPU.scala 52:20]
  reg [31:0] DMemory_892; // @[CPU.scala 52:20]
  reg [31:0] DMemory_893; // @[CPU.scala 52:20]
  reg [31:0] DMemory_894; // @[CPU.scala 52:20]
  reg [31:0] DMemory_895; // @[CPU.scala 52:20]
  reg [31:0] DMemory_896; // @[CPU.scala 52:20]
  reg [31:0] DMemory_897; // @[CPU.scala 52:20]
  reg [31:0] DMemory_898; // @[CPU.scala 52:20]
  reg [31:0] DMemory_899; // @[CPU.scala 52:20]
  reg [31:0] DMemory_900; // @[CPU.scala 52:20]
  reg [31:0] DMemory_901; // @[CPU.scala 52:20]
  reg [31:0] DMemory_902; // @[CPU.scala 52:20]
  reg [31:0] DMemory_903; // @[CPU.scala 52:20]
  reg [31:0] DMemory_904; // @[CPU.scala 52:20]
  reg [31:0] DMemory_905; // @[CPU.scala 52:20]
  reg [31:0] DMemory_906; // @[CPU.scala 52:20]
  reg [31:0] DMemory_907; // @[CPU.scala 52:20]
  reg [31:0] DMemory_908; // @[CPU.scala 52:20]
  reg [31:0] DMemory_909; // @[CPU.scala 52:20]
  reg [31:0] DMemory_910; // @[CPU.scala 52:20]
  reg [31:0] DMemory_911; // @[CPU.scala 52:20]
  reg [31:0] DMemory_912; // @[CPU.scala 52:20]
  reg [31:0] DMemory_913; // @[CPU.scala 52:20]
  reg [31:0] DMemory_914; // @[CPU.scala 52:20]
  reg [31:0] DMemory_915; // @[CPU.scala 52:20]
  reg [31:0] DMemory_916; // @[CPU.scala 52:20]
  reg [31:0] DMemory_917; // @[CPU.scala 52:20]
  reg [31:0] DMemory_918; // @[CPU.scala 52:20]
  reg [31:0] DMemory_919; // @[CPU.scala 52:20]
  reg [31:0] DMemory_920; // @[CPU.scala 52:20]
  reg [31:0] DMemory_921; // @[CPU.scala 52:20]
  reg [31:0] DMemory_922; // @[CPU.scala 52:20]
  reg [31:0] DMemory_923; // @[CPU.scala 52:20]
  reg [31:0] DMemory_924; // @[CPU.scala 52:20]
  reg [31:0] DMemory_925; // @[CPU.scala 52:20]
  reg [31:0] DMemory_926; // @[CPU.scala 52:20]
  reg [31:0] DMemory_927; // @[CPU.scala 52:20]
  reg [31:0] DMemory_928; // @[CPU.scala 52:20]
  reg [31:0] DMemory_929; // @[CPU.scala 52:20]
  reg [31:0] DMemory_930; // @[CPU.scala 52:20]
  reg [31:0] DMemory_931; // @[CPU.scala 52:20]
  reg [31:0] DMemory_932; // @[CPU.scala 52:20]
  reg [31:0] DMemory_933; // @[CPU.scala 52:20]
  reg [31:0] DMemory_934; // @[CPU.scala 52:20]
  reg [31:0] DMemory_935; // @[CPU.scala 52:20]
  reg [31:0] DMemory_936; // @[CPU.scala 52:20]
  reg [31:0] DMemory_937; // @[CPU.scala 52:20]
  reg [31:0] DMemory_938; // @[CPU.scala 52:20]
  reg [31:0] DMemory_939; // @[CPU.scala 52:20]
  reg [31:0] DMemory_940; // @[CPU.scala 52:20]
  reg [31:0] DMemory_941; // @[CPU.scala 52:20]
  reg [31:0] DMemory_942; // @[CPU.scala 52:20]
  reg [31:0] DMemory_943; // @[CPU.scala 52:20]
  reg [31:0] DMemory_944; // @[CPU.scala 52:20]
  reg [31:0] DMemory_945; // @[CPU.scala 52:20]
  reg [31:0] DMemory_946; // @[CPU.scala 52:20]
  reg [31:0] DMemory_947; // @[CPU.scala 52:20]
  reg [31:0] DMemory_948; // @[CPU.scala 52:20]
  reg [31:0] DMemory_949; // @[CPU.scala 52:20]
  reg [31:0] DMemory_950; // @[CPU.scala 52:20]
  reg [31:0] DMemory_951; // @[CPU.scala 52:20]
  reg [31:0] DMemory_952; // @[CPU.scala 52:20]
  reg [31:0] DMemory_953; // @[CPU.scala 52:20]
  reg [31:0] DMemory_954; // @[CPU.scala 52:20]
  reg [31:0] DMemory_955; // @[CPU.scala 52:20]
  reg [31:0] DMemory_956; // @[CPU.scala 52:20]
  reg [31:0] DMemory_957; // @[CPU.scala 52:20]
  reg [31:0] DMemory_958; // @[CPU.scala 52:20]
  reg [31:0] DMemory_959; // @[CPU.scala 52:20]
  reg [31:0] DMemory_960; // @[CPU.scala 52:20]
  reg [31:0] DMemory_961; // @[CPU.scala 52:20]
  reg [31:0] DMemory_962; // @[CPU.scala 52:20]
  reg [31:0] DMemory_963; // @[CPU.scala 52:20]
  reg [31:0] DMemory_964; // @[CPU.scala 52:20]
  reg [31:0] DMemory_965; // @[CPU.scala 52:20]
  reg [31:0] DMemory_966; // @[CPU.scala 52:20]
  reg [31:0] DMemory_967; // @[CPU.scala 52:20]
  reg [31:0] DMemory_968; // @[CPU.scala 52:20]
  reg [31:0] DMemory_969; // @[CPU.scala 52:20]
  reg [31:0] DMemory_970; // @[CPU.scala 52:20]
  reg [31:0] DMemory_971; // @[CPU.scala 52:20]
  reg [31:0] DMemory_972; // @[CPU.scala 52:20]
  reg [31:0] DMemory_973; // @[CPU.scala 52:20]
  reg [31:0] DMemory_974; // @[CPU.scala 52:20]
  reg [31:0] DMemory_975; // @[CPU.scala 52:20]
  reg [31:0] DMemory_976; // @[CPU.scala 52:20]
  reg [31:0] DMemory_977; // @[CPU.scala 52:20]
  reg [31:0] DMemory_978; // @[CPU.scala 52:20]
  reg [31:0] DMemory_979; // @[CPU.scala 52:20]
  reg [31:0] DMemory_980; // @[CPU.scala 52:20]
  reg [31:0] DMemory_981; // @[CPU.scala 52:20]
  reg [31:0] DMemory_982; // @[CPU.scala 52:20]
  reg [31:0] DMemory_983; // @[CPU.scala 52:20]
  reg [31:0] DMemory_984; // @[CPU.scala 52:20]
  reg [31:0] DMemory_985; // @[CPU.scala 52:20]
  reg [31:0] DMemory_986; // @[CPU.scala 52:20]
  reg [31:0] DMemory_987; // @[CPU.scala 52:20]
  reg [31:0] DMemory_988; // @[CPU.scala 52:20]
  reg [31:0] DMemory_989; // @[CPU.scala 52:20]
  reg [31:0] DMemory_990; // @[CPU.scala 52:20]
  reg [31:0] DMemory_991; // @[CPU.scala 52:20]
  reg [31:0] DMemory_992; // @[CPU.scala 52:20]
  reg [31:0] DMemory_993; // @[CPU.scala 52:20]
  reg [31:0] DMemory_994; // @[CPU.scala 52:20]
  reg [31:0] DMemory_995; // @[CPU.scala 52:20]
  reg [31:0] DMemory_996; // @[CPU.scala 52:20]
  reg [31:0] DMemory_997; // @[CPU.scala 52:20]
  reg [31:0] DMemory_998; // @[CPU.scala 52:20]
  reg [31:0] DMemory_999; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1000; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1001; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1002; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1003; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1004; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1005; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1006; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1007; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1008; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1009; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1010; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1011; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1012; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1013; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1014; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1015; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1016; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1017; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1018; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1019; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1020; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1021; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1022; // @[CPU.scala 52:20]
  reg [31:0] DMemory_1023; // @[CPU.scala 52:20]
  reg [31:0] IMemory_0; // @[CPU.scala 53:20]
  reg [31:0] IMemory_1; // @[CPU.scala 53:20]
  reg [31:0] IMemory_2; // @[CPU.scala 53:20]
  reg [31:0] IMemory_3; // @[CPU.scala 53:20]
  reg [31:0] IFIDIR; // @[CPU.scala 54:49]
  reg [31:0] IDEXIR; // @[CPU.scala 54:49]
  reg [31:0] EXMEMIR; // @[CPU.scala 54:49]
  reg [31:0] MEMWBIR; // @[CPU.scala 54:49]
  reg [63:0] CurPC; // @[CPU.scala 57:22]
  wire [4:0] EXMEMrd = EXMEMIR[11:7]; // @[CPU.scala 89:32]
  wire [4:0] IDEXrd = IDEXIR[11:7]; // @[CPU.scala 90:30]
  wire [2:0] IFID_funct3 = IFIDIR[14:12]; // @[CPU.scala 91:29]
  wire [4:0] IFIDrs1 = io_rvfi_rst ? IFIDIR[19:15] : IFIDIR[19:15]; // @[CPU.scala 61:21 64:13 81:13]
  wire [4:0] MEMWBrd = io_rvfi_rst ? MEMWBIR[11:7] : MEMWBIR[11:7]; // @[CPU.scala 61:21 70:13 87:13]
  wire  _bypassAFromWB_T_1 = IFIDrs1 != 5'h0; // @[CPU.scala 94:41]
  wire [6:0] MEMWBop = io_rvfi_rst ? MEMWBIR[6:0] : MEMWBIR[6:0]; // @[CPU.scala 61:21 69:13 86:13]
  wire  _bypassAFromWB_T_3 = MEMWBop == 7'h33; // @[CPU.scala 94:62]
  wire  _bypassAFromWB_T_4 = MEMWBop == 7'h3; // @[CPU.scala 94:83]
  wire  _bypassAFromWB_T_5 = MEMWBop == 7'h33 | MEMWBop == 7'h3; // @[CPU.scala 94:72]
  wire  bypassAFromWB = IFIDrs1 == MEMWBrd & IFIDrs1 != 5'h0 & (MEMWBop == 7'h33 | MEMWBop == 7'h3); // @[CPU.scala 94:50]
  wire [4:0] IFIDrs2 = io_rvfi_rst ? IFIDIR[24:20] : IFIDIR[24:20]; // @[CPU.scala 61:21 65:13 82:13]
  wire  _bypassBFromWB_T_1 = IFIDrs2 != 5'h0; // @[CPU.scala 96:41]
  wire  bypassBFromWB = IFIDrs2 == MEMWBrd & IFIDrs2 != 5'h0 & _bypassAFromWB_T_5; // @[CPU.scala 96:50]
  wire  _bypassAFromMEM_T_2 = IFIDrs1 == EXMEMrd & _bypassAFromWB_T_1; // @[CPU.scala 98:29]
  wire [6:0] EXMEMop = io_rvfi_rst ? EXMEMIR[6:0] : EXMEMIR[6:0]; // @[CPU.scala 61:21 68:13 85:13]
  wire  _bypassAFromMEM_T_3 = EXMEMop == 7'h33; // @[CPU.scala 98:62]
  wire  bypassAFromMEM = IFIDrs1 == EXMEMrd & _bypassAFromWB_T_1 & EXMEMop == 7'h33; // @[CPU.scala 98:50]
  wire  _bypassBFromMEM_T_2 = IFIDrs2 == EXMEMrd & _bypassBFromWB_T_1; // @[CPU.scala 100:29]
  wire  bypassBFromMEM = IFIDrs2 == EXMEMrd & _bypassBFromWB_T_1 & _bypassAFromMEM_T_3; // @[CPU.scala 100:50]
  wire  _bypassAFromEX_T_2 = IFIDrs1 == IDEXrd & _bypassAFromWB_T_1; // @[CPU.scala 102:28]
  wire [6:0] IDEXop = io_rvfi_rst ? IDEXIR[6:0] : IDEXIR[6:0]; // @[CPU.scala 61:21 66:12 83:12]
  wire  _bypassAFromEX_T_3 = IDEXop == 7'h33; // @[CPU.scala 102:60]
  wire  bypassAFromEX = IFIDrs1 == IDEXrd & _bypassAFromWB_T_1 & IDEXop == 7'h33; // @[CPU.scala 102:49]
  wire  _bypassBFromEX_T_2 = IFIDrs2 == IDEXrd & _bypassBFromWB_T_1; // @[CPU.scala 104:28]
  wire  bypassBFromEX = IFIDrs2 == IDEXrd & _bypassBFromWB_T_1 & _bypassAFromEX_T_3; // @[CPU.scala 104:49]
  wire  _stall_T = EXMEMop == 7'h3; // @[CPU.scala 107:16]
  wire  _stall_T_8 = EXMEMop == 7'h3 & (_bypassAFromMEM_T_2 | _bypassBFromMEM_T_2); // @[CPU.scala 107:24]
  wire  _stall_T_9 = IDEXop == 7'h3; // @[CPU.scala 109:15]
  wire  _stall_T_17 = IDEXop == 7'h3 & (_bypassAFromEX_T_2 | _bypassBFromEX_T_2); // @[CPU.scala 109:23]
  wire  stall = _stall_T_8 | _stall_T_17; // @[CPU.scala 108:7]
  wire [6:0] IFIDop = io_rvfi_rst ? IFIDIR[6:0] : IFIDIR[6:0]; // @[CPU.scala 61:21 67:12 84:12]
  wire [63:0] _A_T_1 = IDEXA + IDEXB; // @[CPU.scala 150:20]
  wire [63:0] _GEN_3141 = 5'h1 == IFIDrs1 ? Regs_1 : Regs_0; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3142 = 5'h2 == IFIDrs1 ? Regs_2 : _GEN_3141; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3143 = 5'h3 == IFIDrs1 ? Regs_3 : _GEN_3142; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3144 = 5'h4 == IFIDrs1 ? Regs_4 : _GEN_3143; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3145 = 5'h5 == IFIDrs1 ? Regs_5 : _GEN_3144; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3146 = 5'h6 == IFIDrs1 ? Regs_6 : _GEN_3145; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3147 = 5'h7 == IFIDrs1 ? Regs_7 : _GEN_3146; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3148 = 5'h8 == IFIDrs1 ? Regs_8 : _GEN_3147; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3149 = 5'h9 == IFIDrs1 ? Regs_9 : _GEN_3148; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3150 = 5'ha == IFIDrs1 ? Regs_10 : _GEN_3149; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3151 = 5'hb == IFIDrs1 ? Regs_11 : _GEN_3150; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3152 = 5'hc == IFIDrs1 ? Regs_12 : _GEN_3151; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3153 = 5'hd == IFIDrs1 ? Regs_13 : _GEN_3152; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3154 = 5'he == IFIDrs1 ? Regs_14 : _GEN_3153; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3155 = 5'hf == IFIDrs1 ? Regs_15 : _GEN_3154; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3156 = 5'h10 == IFIDrs1 ? Regs_16 : _GEN_3155; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3157 = 5'h11 == IFIDrs1 ? Regs_17 : _GEN_3156; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3158 = 5'h12 == IFIDrs1 ? Regs_18 : _GEN_3157; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3159 = 5'h13 == IFIDrs1 ? Regs_19 : _GEN_3158; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3160 = 5'h14 == IFIDrs1 ? Regs_20 : _GEN_3159; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3161 = 5'h15 == IFIDrs1 ? Regs_21 : _GEN_3160; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3162 = 5'h16 == IFIDrs1 ? Regs_22 : _GEN_3161; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3163 = 5'h17 == IFIDrs1 ? Regs_23 : _GEN_3162; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3164 = 5'h18 == IFIDrs1 ? Regs_24 : _GEN_3163; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3165 = 5'h19 == IFIDrs1 ? Regs_25 : _GEN_3164; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3166 = 5'h1a == IFIDrs1 ? Regs_26 : _GEN_3165; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3167 = 5'h1b == IFIDrs1 ? Regs_27 : _GEN_3166; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3168 = 5'h1c == IFIDrs1 ? Regs_28 : _GEN_3167; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3169 = 5'h1d == IFIDrs1 ? Regs_29 : _GEN_3168; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3170 = 5'h1e == IFIDrs1 ? Regs_30 : _GEN_3169; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3171 = 5'h1f == IFIDrs1 ? Regs_31 : _GEN_3170; // @[CPU.scala 158:{15,15}]
  wire [63:0] _GEN_3173 = bypassAFromWB ? MEMWBValue : _GEN_3171; // @[CPU.scala 154:33 156:11 159:11]
  wire [63:0] _GEN_3175 = bypassAFromMEM ? EXMEMALUOut : _GEN_3173; // @[CPU.scala 151:34 153:11]
  wire [63:0] _GEN_3177 = bypassAFromEX ? _A_T_1 : _GEN_3175; // @[CPU.scala 148:27 150:11]
  wire [63:0] A = ~stall ? _GEN_3177 : 64'h0; // @[CPU.scala 121:27]
  wire [63:0] _B_T_1 = IDEXB + IDEXA; // @[CPU.scala 163:20]
  wire [63:0] _GEN_3179 = 5'h1 == IFIDrs2 ? Regs_1 : Regs_0; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3180 = 5'h2 == IFIDrs2 ? Regs_2 : _GEN_3179; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3181 = 5'h3 == IFIDrs2 ? Regs_3 : _GEN_3180; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3182 = 5'h4 == IFIDrs2 ? Regs_4 : _GEN_3181; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3183 = 5'h5 == IFIDrs2 ? Regs_5 : _GEN_3182; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3184 = 5'h6 == IFIDrs2 ? Regs_6 : _GEN_3183; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3185 = 5'h7 == IFIDrs2 ? Regs_7 : _GEN_3184; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3186 = 5'h8 == IFIDrs2 ? Regs_8 : _GEN_3185; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3187 = 5'h9 == IFIDrs2 ? Regs_9 : _GEN_3186; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3188 = 5'ha == IFIDrs2 ? Regs_10 : _GEN_3187; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3189 = 5'hb == IFIDrs2 ? Regs_11 : _GEN_3188; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3190 = 5'hc == IFIDrs2 ? Regs_12 : _GEN_3189; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3191 = 5'hd == IFIDrs2 ? Regs_13 : _GEN_3190; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3192 = 5'he == IFIDrs2 ? Regs_14 : _GEN_3191; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3193 = 5'hf == IFIDrs2 ? Regs_15 : _GEN_3192; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3194 = 5'h10 == IFIDrs2 ? Regs_16 : _GEN_3193; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3195 = 5'h11 == IFIDrs2 ? Regs_17 : _GEN_3194; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3196 = 5'h12 == IFIDrs2 ? Regs_18 : _GEN_3195; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3197 = 5'h13 == IFIDrs2 ? Regs_19 : _GEN_3196; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3198 = 5'h14 == IFIDrs2 ? Regs_20 : _GEN_3197; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3199 = 5'h15 == IFIDrs2 ? Regs_21 : _GEN_3198; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3200 = 5'h16 == IFIDrs2 ? Regs_22 : _GEN_3199; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3201 = 5'h17 == IFIDrs2 ? Regs_23 : _GEN_3200; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3202 = 5'h18 == IFIDrs2 ? Regs_24 : _GEN_3201; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3203 = 5'h19 == IFIDrs2 ? Regs_25 : _GEN_3202; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3204 = 5'h1a == IFIDrs2 ? Regs_26 : _GEN_3203; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3205 = 5'h1b == IFIDrs2 ? Regs_27 : _GEN_3204; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3206 = 5'h1c == IFIDrs2 ? Regs_28 : _GEN_3205; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3207 = 5'h1d == IFIDrs2 ? Regs_29 : _GEN_3206; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3208 = 5'h1e == IFIDrs2 ? Regs_30 : _GEN_3207; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3209 = 5'h1f == IFIDrs2 ? Regs_31 : _GEN_3208; // @[CPU.scala 171:{15,15}]
  wire [63:0] _GEN_3211 = bypassBFromWB ? MEMWBValue : _GEN_3209; // @[CPU.scala 167:33 169:11 172:11]
  wire [63:0] _GEN_3213 = bypassBFromMEM ? EXMEMALUOut : _GEN_3211; // @[CPU.scala 164:34 166:11]
  wire [63:0] _GEN_3215 = bypassBFromEX ? _B_T_1 : _GEN_3213; // @[CPU.scala 161:27 163:11]
  wire [63:0] B = ~stall ? _GEN_3215 : 64'h0; // @[CPU.scala 121:27]
  wire  takeBranch = IFIDop == 7'h63 & IFID_funct3 == 3'h0 & A == B; // @[CPU.scala 113:64]
  wire [63:0] _IFIDIR_T = {{2'd0}, PC[63:2]}; // @[CPU.scala 125:31]
  wire [31:0] _GEN_2113 = 10'h1 == _IFIDIR_T[9:0] ? IMemory_1 : IMemory_0; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2114 = 10'h2 == _IFIDIR_T[9:0] ? IMemory_2 : _GEN_2113; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2115 = 10'h3 == _IFIDIR_T[9:0] ? IMemory_3 : _GEN_2114; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2116 = 10'h4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2115; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2117 = 10'h5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2116; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2118 = 10'h6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2117; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2119 = 10'h7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2118; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2120 = 10'h8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2119; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2121 = 10'h9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2120; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2122 = 10'ha == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2121; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2123 = 10'hb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2122; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2124 = 10'hc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2123; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2125 = 10'hd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2124; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2126 = 10'he == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2125; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2127 = 10'hf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2126; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2128 = 10'h10 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2127; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2129 = 10'h11 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2128; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2130 = 10'h12 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2129; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2131 = 10'h13 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2130; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2132 = 10'h14 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2131; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2133 = 10'h15 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2132; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2134 = 10'h16 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2133; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2135 = 10'h17 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2134; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2136 = 10'h18 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2135; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2137 = 10'h19 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2136; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2138 = 10'h1a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2137; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2139 = 10'h1b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2138; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2140 = 10'h1c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2139; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2141 = 10'h1d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2140; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2142 = 10'h1e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2141; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2143 = 10'h1f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2142; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2144 = 10'h20 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2143; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2145 = 10'h21 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2144; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2146 = 10'h22 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2145; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2147 = 10'h23 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2146; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2148 = 10'h24 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2147; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2149 = 10'h25 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2148; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2150 = 10'h26 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2149; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2151 = 10'h27 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2150; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2152 = 10'h28 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2151; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2153 = 10'h29 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2152; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2154 = 10'h2a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2153; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2155 = 10'h2b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2154; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2156 = 10'h2c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2155; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2157 = 10'h2d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2156; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2158 = 10'h2e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2157; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2159 = 10'h2f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2158; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2160 = 10'h30 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2159; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2161 = 10'h31 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2160; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2162 = 10'h32 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2161; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2163 = 10'h33 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2162; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2164 = 10'h34 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2163; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2165 = 10'h35 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2164; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2166 = 10'h36 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2165; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2167 = 10'h37 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2166; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2168 = 10'h38 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2167; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2169 = 10'h39 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2168; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2170 = 10'h3a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2169; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2171 = 10'h3b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2170; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2172 = 10'h3c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2171; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2173 = 10'h3d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2172; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2174 = 10'h3e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2173; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2175 = 10'h3f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2174; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2176 = 10'h40 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2175; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2177 = 10'h41 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2176; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2178 = 10'h42 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2177; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2179 = 10'h43 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2178; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2180 = 10'h44 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2179; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2181 = 10'h45 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2180; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2182 = 10'h46 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2181; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2183 = 10'h47 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2182; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2184 = 10'h48 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2183; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2185 = 10'h49 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2184; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2186 = 10'h4a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2185; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2187 = 10'h4b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2186; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2188 = 10'h4c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2187; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2189 = 10'h4d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2188; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2190 = 10'h4e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2189; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2191 = 10'h4f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2190; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2192 = 10'h50 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2191; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2193 = 10'h51 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2192; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2194 = 10'h52 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2193; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2195 = 10'h53 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2194; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2196 = 10'h54 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2195; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2197 = 10'h55 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2196; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2198 = 10'h56 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2197; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2199 = 10'h57 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2198; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2200 = 10'h58 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2199; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2201 = 10'h59 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2200; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2202 = 10'h5a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2201; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2203 = 10'h5b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2202; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2204 = 10'h5c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2203; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2205 = 10'h5d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2204; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2206 = 10'h5e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2205; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2207 = 10'h5f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2206; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2208 = 10'h60 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2207; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2209 = 10'h61 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2208; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2210 = 10'h62 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2209; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2211 = 10'h63 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2210; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2212 = 10'h64 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2211; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2213 = 10'h65 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2212; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2214 = 10'h66 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2213; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2215 = 10'h67 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2214; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2216 = 10'h68 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2215; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2217 = 10'h69 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2216; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2218 = 10'h6a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2217; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2219 = 10'h6b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2218; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2220 = 10'h6c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2219; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2221 = 10'h6d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2220; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2222 = 10'h6e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2221; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2223 = 10'h6f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2222; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2224 = 10'h70 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2223; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2225 = 10'h71 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2224; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2226 = 10'h72 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2225; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2227 = 10'h73 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2226; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2228 = 10'h74 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2227; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2229 = 10'h75 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2228; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2230 = 10'h76 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2229; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2231 = 10'h77 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2230; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2232 = 10'h78 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2231; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2233 = 10'h79 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2232; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2234 = 10'h7a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2233; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2235 = 10'h7b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2234; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2236 = 10'h7c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2235; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2237 = 10'h7d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2236; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2238 = 10'h7e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2237; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2239 = 10'h7f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2238; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2240 = 10'h80 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2239; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2241 = 10'h81 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2240; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2242 = 10'h82 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2241; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2243 = 10'h83 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2242; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2244 = 10'h84 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2243; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2245 = 10'h85 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2244; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2246 = 10'h86 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2245; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2247 = 10'h87 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2246; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2248 = 10'h88 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2247; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2249 = 10'h89 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2248; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2250 = 10'h8a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2249; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2251 = 10'h8b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2250; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2252 = 10'h8c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2251; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2253 = 10'h8d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2252; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2254 = 10'h8e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2253; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2255 = 10'h8f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2254; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2256 = 10'h90 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2255; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2257 = 10'h91 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2256; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2258 = 10'h92 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2257; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2259 = 10'h93 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2258; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2260 = 10'h94 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2259; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2261 = 10'h95 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2260; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2262 = 10'h96 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2261; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2263 = 10'h97 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2262; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2264 = 10'h98 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2263; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2265 = 10'h99 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2264; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2266 = 10'h9a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2265; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2267 = 10'h9b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2266; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2268 = 10'h9c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2267; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2269 = 10'h9d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2268; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2270 = 10'h9e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2269; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2271 = 10'h9f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2270; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2272 = 10'ha0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2271; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2273 = 10'ha1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2272; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2274 = 10'ha2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2273; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2275 = 10'ha3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2274; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2276 = 10'ha4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2275; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2277 = 10'ha5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2276; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2278 = 10'ha6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2277; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2279 = 10'ha7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2278; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2280 = 10'ha8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2279; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2281 = 10'ha9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2280; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2282 = 10'haa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2281; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2283 = 10'hab == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2282; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2284 = 10'hac == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2283; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2285 = 10'had == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2284; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2286 = 10'hae == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2285; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2287 = 10'haf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2286; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2288 = 10'hb0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2287; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2289 = 10'hb1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2288; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2290 = 10'hb2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2289; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2291 = 10'hb3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2290; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2292 = 10'hb4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2291; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2293 = 10'hb5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2292; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2294 = 10'hb6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2293; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2295 = 10'hb7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2294; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2296 = 10'hb8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2295; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2297 = 10'hb9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2296; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2298 = 10'hba == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2297; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2299 = 10'hbb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2298; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2300 = 10'hbc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2299; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2301 = 10'hbd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2300; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2302 = 10'hbe == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2301; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2303 = 10'hbf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2302; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2304 = 10'hc0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2303; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2305 = 10'hc1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2304; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2306 = 10'hc2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2305; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2307 = 10'hc3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2306; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2308 = 10'hc4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2307; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2309 = 10'hc5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2308; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2310 = 10'hc6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2309; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2311 = 10'hc7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2310; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2312 = 10'hc8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2311; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2313 = 10'hc9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2312; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2314 = 10'hca == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2313; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2315 = 10'hcb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2314; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2316 = 10'hcc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2315; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2317 = 10'hcd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2316; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2318 = 10'hce == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2317; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2319 = 10'hcf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2318; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2320 = 10'hd0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2319; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2321 = 10'hd1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2320; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2322 = 10'hd2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2321; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2323 = 10'hd3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2322; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2324 = 10'hd4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2323; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2325 = 10'hd5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2324; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2326 = 10'hd6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2325; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2327 = 10'hd7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2326; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2328 = 10'hd8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2327; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2329 = 10'hd9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2328; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2330 = 10'hda == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2329; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2331 = 10'hdb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2330; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2332 = 10'hdc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2331; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2333 = 10'hdd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2332; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2334 = 10'hde == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2333; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2335 = 10'hdf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2334; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2336 = 10'he0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2335; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2337 = 10'he1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2336; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2338 = 10'he2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2337; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2339 = 10'he3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2338; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2340 = 10'he4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2339; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2341 = 10'he5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2340; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2342 = 10'he6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2341; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2343 = 10'he7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2342; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2344 = 10'he8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2343; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2345 = 10'he9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2344; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2346 = 10'hea == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2345; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2347 = 10'heb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2346; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2348 = 10'hec == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2347; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2349 = 10'hed == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2348; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2350 = 10'hee == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2349; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2351 = 10'hef == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2350; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2352 = 10'hf0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2351; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2353 = 10'hf1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2352; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2354 = 10'hf2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2353; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2355 = 10'hf3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2354; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2356 = 10'hf4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2355; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2357 = 10'hf5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2356; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2358 = 10'hf6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2357; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2359 = 10'hf7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2358; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2360 = 10'hf8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2359; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2361 = 10'hf9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2360; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2362 = 10'hfa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2361; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2363 = 10'hfb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2362; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2364 = 10'hfc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2363; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2365 = 10'hfd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2364; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2366 = 10'hfe == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2365; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2367 = 10'hff == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2366; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2368 = 10'h100 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2367; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2369 = 10'h101 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2368; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2370 = 10'h102 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2369; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2371 = 10'h103 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2370; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2372 = 10'h104 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2371; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2373 = 10'h105 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2372; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2374 = 10'h106 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2373; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2375 = 10'h107 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2374; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2376 = 10'h108 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2375; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2377 = 10'h109 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2376; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2378 = 10'h10a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2377; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2379 = 10'h10b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2378; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2380 = 10'h10c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2379; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2381 = 10'h10d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2380; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2382 = 10'h10e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2381; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2383 = 10'h10f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2382; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2384 = 10'h110 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2383; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2385 = 10'h111 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2384; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2386 = 10'h112 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2385; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2387 = 10'h113 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2386; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2388 = 10'h114 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2387; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2389 = 10'h115 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2388; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2390 = 10'h116 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2389; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2391 = 10'h117 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2390; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2392 = 10'h118 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2391; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2393 = 10'h119 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2392; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2394 = 10'h11a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2393; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2395 = 10'h11b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2394; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2396 = 10'h11c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2395; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2397 = 10'h11d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2396; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2398 = 10'h11e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2397; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2399 = 10'h11f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2398; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2400 = 10'h120 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2399; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2401 = 10'h121 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2400; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2402 = 10'h122 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2401; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2403 = 10'h123 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2402; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2404 = 10'h124 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2403; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2405 = 10'h125 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2404; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2406 = 10'h126 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2405; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2407 = 10'h127 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2406; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2408 = 10'h128 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2407; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2409 = 10'h129 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2408; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2410 = 10'h12a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2409; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2411 = 10'h12b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2410; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2412 = 10'h12c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2411; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2413 = 10'h12d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2412; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2414 = 10'h12e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2413; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2415 = 10'h12f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2414; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2416 = 10'h130 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2415; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2417 = 10'h131 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2416; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2418 = 10'h132 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2417; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2419 = 10'h133 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2418; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2420 = 10'h134 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2419; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2421 = 10'h135 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2420; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2422 = 10'h136 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2421; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2423 = 10'h137 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2422; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2424 = 10'h138 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2423; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2425 = 10'h139 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2424; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2426 = 10'h13a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2425; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2427 = 10'h13b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2426; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2428 = 10'h13c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2427; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2429 = 10'h13d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2428; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2430 = 10'h13e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2429; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2431 = 10'h13f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2430; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2432 = 10'h140 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2431; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2433 = 10'h141 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2432; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2434 = 10'h142 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2433; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2435 = 10'h143 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2434; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2436 = 10'h144 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2435; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2437 = 10'h145 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2436; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2438 = 10'h146 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2437; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2439 = 10'h147 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2438; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2440 = 10'h148 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2439; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2441 = 10'h149 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2440; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2442 = 10'h14a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2441; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2443 = 10'h14b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2442; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2444 = 10'h14c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2443; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2445 = 10'h14d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2444; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2446 = 10'h14e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2445; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2447 = 10'h14f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2446; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2448 = 10'h150 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2447; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2449 = 10'h151 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2448; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2450 = 10'h152 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2449; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2451 = 10'h153 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2450; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2452 = 10'h154 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2451; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2453 = 10'h155 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2452; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2454 = 10'h156 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2453; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2455 = 10'h157 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2454; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2456 = 10'h158 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2455; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2457 = 10'h159 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2456; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2458 = 10'h15a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2457; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2459 = 10'h15b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2458; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2460 = 10'h15c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2459; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2461 = 10'h15d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2460; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2462 = 10'h15e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2461; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2463 = 10'h15f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2462; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2464 = 10'h160 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2463; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2465 = 10'h161 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2464; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2466 = 10'h162 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2465; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2467 = 10'h163 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2466; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2468 = 10'h164 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2467; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2469 = 10'h165 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2468; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2470 = 10'h166 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2469; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2471 = 10'h167 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2470; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2472 = 10'h168 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2471; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2473 = 10'h169 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2472; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2474 = 10'h16a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2473; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2475 = 10'h16b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2474; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2476 = 10'h16c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2475; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2477 = 10'h16d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2476; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2478 = 10'h16e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2477; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2479 = 10'h16f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2478; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2480 = 10'h170 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2479; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2481 = 10'h171 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2480; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2482 = 10'h172 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2481; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2483 = 10'h173 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2482; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2484 = 10'h174 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2483; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2485 = 10'h175 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2484; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2486 = 10'h176 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2485; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2487 = 10'h177 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2486; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2488 = 10'h178 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2487; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2489 = 10'h179 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2488; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2490 = 10'h17a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2489; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2491 = 10'h17b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2490; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2492 = 10'h17c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2491; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2493 = 10'h17d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2492; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2494 = 10'h17e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2493; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2495 = 10'h17f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2494; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2496 = 10'h180 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2495; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2497 = 10'h181 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2496; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2498 = 10'h182 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2497; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2499 = 10'h183 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2498; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2500 = 10'h184 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2499; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2501 = 10'h185 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2500; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2502 = 10'h186 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2501; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2503 = 10'h187 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2502; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2504 = 10'h188 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2503; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2505 = 10'h189 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2504; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2506 = 10'h18a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2505; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2507 = 10'h18b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2506; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2508 = 10'h18c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2507; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2509 = 10'h18d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2508; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2510 = 10'h18e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2509; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2511 = 10'h18f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2510; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2512 = 10'h190 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2511; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2513 = 10'h191 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2512; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2514 = 10'h192 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2513; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2515 = 10'h193 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2514; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2516 = 10'h194 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2515; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2517 = 10'h195 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2516; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2518 = 10'h196 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2517; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2519 = 10'h197 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2518; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2520 = 10'h198 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2519; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2521 = 10'h199 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2520; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2522 = 10'h19a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2521; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2523 = 10'h19b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2522; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2524 = 10'h19c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2523; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2525 = 10'h19d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2524; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2526 = 10'h19e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2525; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2527 = 10'h19f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2526; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2528 = 10'h1a0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2527; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2529 = 10'h1a1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2528; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2530 = 10'h1a2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2529; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2531 = 10'h1a3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2530; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2532 = 10'h1a4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2531; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2533 = 10'h1a5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2532; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2534 = 10'h1a6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2533; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2535 = 10'h1a7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2534; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2536 = 10'h1a8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2535; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2537 = 10'h1a9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2536; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2538 = 10'h1aa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2537; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2539 = 10'h1ab == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2538; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2540 = 10'h1ac == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2539; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2541 = 10'h1ad == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2540; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2542 = 10'h1ae == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2541; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2543 = 10'h1af == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2542; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2544 = 10'h1b0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2543; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2545 = 10'h1b1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2544; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2546 = 10'h1b2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2545; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2547 = 10'h1b3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2546; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2548 = 10'h1b4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2547; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2549 = 10'h1b5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2548; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2550 = 10'h1b6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2549; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2551 = 10'h1b7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2550; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2552 = 10'h1b8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2551; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2553 = 10'h1b9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2552; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2554 = 10'h1ba == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2553; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2555 = 10'h1bb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2554; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2556 = 10'h1bc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2555; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2557 = 10'h1bd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2556; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2558 = 10'h1be == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2557; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2559 = 10'h1bf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2558; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2560 = 10'h1c0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2559; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2561 = 10'h1c1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2560; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2562 = 10'h1c2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2561; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2563 = 10'h1c3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2562; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2564 = 10'h1c4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2563; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2565 = 10'h1c5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2564; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2566 = 10'h1c6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2565; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2567 = 10'h1c7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2566; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2568 = 10'h1c8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2567; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2569 = 10'h1c9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2568; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2570 = 10'h1ca == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2569; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2571 = 10'h1cb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2570; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2572 = 10'h1cc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2571; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2573 = 10'h1cd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2572; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2574 = 10'h1ce == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2573; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2575 = 10'h1cf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2574; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2576 = 10'h1d0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2575; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2577 = 10'h1d1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2576; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2578 = 10'h1d2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2577; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2579 = 10'h1d3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2578; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2580 = 10'h1d4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2579; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2581 = 10'h1d5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2580; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2582 = 10'h1d6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2581; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2583 = 10'h1d7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2582; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2584 = 10'h1d8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2583; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2585 = 10'h1d9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2584; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2586 = 10'h1da == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2585; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2587 = 10'h1db == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2586; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2588 = 10'h1dc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2587; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2589 = 10'h1dd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2588; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2590 = 10'h1de == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2589; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2591 = 10'h1df == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2590; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2592 = 10'h1e0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2591; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2593 = 10'h1e1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2592; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2594 = 10'h1e2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2593; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2595 = 10'h1e3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2594; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2596 = 10'h1e4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2595; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2597 = 10'h1e5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2596; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2598 = 10'h1e6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2597; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2599 = 10'h1e7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2598; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2600 = 10'h1e8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2599; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2601 = 10'h1e9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2600; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2602 = 10'h1ea == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2601; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2603 = 10'h1eb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2602; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2604 = 10'h1ec == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2603; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2605 = 10'h1ed == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2604; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2606 = 10'h1ee == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2605; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2607 = 10'h1ef == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2606; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2608 = 10'h1f0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2607; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2609 = 10'h1f1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2608; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2610 = 10'h1f2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2609; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2611 = 10'h1f3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2610; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2612 = 10'h1f4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2611; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2613 = 10'h1f5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2612; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2614 = 10'h1f6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2613; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2615 = 10'h1f7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2614; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2616 = 10'h1f8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2615; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2617 = 10'h1f9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2616; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2618 = 10'h1fa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2617; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2619 = 10'h1fb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2618; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2620 = 10'h1fc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2619; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2621 = 10'h1fd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2620; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2622 = 10'h1fe == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2621; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2623 = 10'h1ff == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2622; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2624 = 10'h200 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2623; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2625 = 10'h201 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2624; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2626 = 10'h202 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2625; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2627 = 10'h203 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2626; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2628 = 10'h204 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2627; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2629 = 10'h205 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2628; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2630 = 10'h206 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2629; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2631 = 10'h207 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2630; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2632 = 10'h208 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2631; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2633 = 10'h209 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2632; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2634 = 10'h20a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2633; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2635 = 10'h20b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2634; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2636 = 10'h20c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2635; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2637 = 10'h20d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2636; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2638 = 10'h20e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2637; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2639 = 10'h20f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2638; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2640 = 10'h210 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2639; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2641 = 10'h211 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2640; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2642 = 10'h212 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2641; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2643 = 10'h213 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2642; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2644 = 10'h214 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2643; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2645 = 10'h215 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2644; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2646 = 10'h216 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2645; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2647 = 10'h217 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2646; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2648 = 10'h218 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2647; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2649 = 10'h219 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2648; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2650 = 10'h21a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2649; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2651 = 10'h21b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2650; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2652 = 10'h21c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2651; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2653 = 10'h21d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2652; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2654 = 10'h21e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2653; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2655 = 10'h21f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2654; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2656 = 10'h220 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2655; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2657 = 10'h221 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2656; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2658 = 10'h222 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2657; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2659 = 10'h223 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2658; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2660 = 10'h224 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2659; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2661 = 10'h225 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2660; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2662 = 10'h226 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2661; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2663 = 10'h227 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2662; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2664 = 10'h228 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2663; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2665 = 10'h229 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2664; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2666 = 10'h22a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2665; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2667 = 10'h22b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2666; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2668 = 10'h22c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2667; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2669 = 10'h22d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2668; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2670 = 10'h22e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2669; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2671 = 10'h22f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2670; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2672 = 10'h230 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2671; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2673 = 10'h231 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2672; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2674 = 10'h232 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2673; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2675 = 10'h233 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2674; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2676 = 10'h234 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2675; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2677 = 10'h235 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2676; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2678 = 10'h236 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2677; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2679 = 10'h237 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2678; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2680 = 10'h238 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2679; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2681 = 10'h239 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2680; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2682 = 10'h23a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2681; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2683 = 10'h23b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2682; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2684 = 10'h23c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2683; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2685 = 10'h23d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2684; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2686 = 10'h23e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2685; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2687 = 10'h23f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2686; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2688 = 10'h240 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2687; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2689 = 10'h241 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2688; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2690 = 10'h242 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2689; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2691 = 10'h243 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2690; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2692 = 10'h244 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2691; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2693 = 10'h245 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2692; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2694 = 10'h246 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2693; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2695 = 10'h247 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2694; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2696 = 10'h248 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2695; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2697 = 10'h249 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2696; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2698 = 10'h24a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2697; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2699 = 10'h24b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2698; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2700 = 10'h24c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2699; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2701 = 10'h24d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2700; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2702 = 10'h24e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2701; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2703 = 10'h24f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2702; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2704 = 10'h250 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2703; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2705 = 10'h251 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2704; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2706 = 10'h252 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2705; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2707 = 10'h253 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2706; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2708 = 10'h254 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2707; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2709 = 10'h255 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2708; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2710 = 10'h256 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2709; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2711 = 10'h257 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2710; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2712 = 10'h258 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2711; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2713 = 10'h259 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2712; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2714 = 10'h25a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2713; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2715 = 10'h25b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2714; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2716 = 10'h25c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2715; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2717 = 10'h25d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2716; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2718 = 10'h25e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2717; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2719 = 10'h25f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2718; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2720 = 10'h260 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2719; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2721 = 10'h261 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2720; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2722 = 10'h262 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2721; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2723 = 10'h263 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2722; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2724 = 10'h264 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2723; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2725 = 10'h265 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2724; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2726 = 10'h266 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2725; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2727 = 10'h267 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2726; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2728 = 10'h268 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2727; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2729 = 10'h269 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2728; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2730 = 10'h26a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2729; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2731 = 10'h26b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2730; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2732 = 10'h26c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2731; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2733 = 10'h26d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2732; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2734 = 10'h26e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2733; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2735 = 10'h26f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2734; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2736 = 10'h270 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2735; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2737 = 10'h271 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2736; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2738 = 10'h272 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2737; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2739 = 10'h273 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2738; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2740 = 10'h274 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2739; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2741 = 10'h275 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2740; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2742 = 10'h276 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2741; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2743 = 10'h277 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2742; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2744 = 10'h278 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2743; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2745 = 10'h279 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2744; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2746 = 10'h27a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2745; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2747 = 10'h27b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2746; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2748 = 10'h27c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2747; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2749 = 10'h27d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2748; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2750 = 10'h27e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2749; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2751 = 10'h27f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2750; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2752 = 10'h280 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2751; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2753 = 10'h281 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2752; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2754 = 10'h282 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2753; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2755 = 10'h283 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2754; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2756 = 10'h284 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2755; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2757 = 10'h285 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2756; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2758 = 10'h286 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2757; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2759 = 10'h287 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2758; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2760 = 10'h288 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2759; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2761 = 10'h289 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2760; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2762 = 10'h28a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2761; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2763 = 10'h28b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2762; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2764 = 10'h28c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2763; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2765 = 10'h28d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2764; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2766 = 10'h28e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2765; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2767 = 10'h28f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2766; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2768 = 10'h290 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2767; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2769 = 10'h291 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2768; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2770 = 10'h292 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2769; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2771 = 10'h293 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2770; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2772 = 10'h294 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2771; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2773 = 10'h295 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2772; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2774 = 10'h296 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2773; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2775 = 10'h297 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2774; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2776 = 10'h298 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2775; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2777 = 10'h299 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2776; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2778 = 10'h29a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2777; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2779 = 10'h29b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2778; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2780 = 10'h29c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2779; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2781 = 10'h29d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2780; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2782 = 10'h29e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2781; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2783 = 10'h29f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2782; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2784 = 10'h2a0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2783; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2785 = 10'h2a1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2784; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2786 = 10'h2a2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2785; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2787 = 10'h2a3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2786; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2788 = 10'h2a4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2787; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2789 = 10'h2a5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2788; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2790 = 10'h2a6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2789; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2791 = 10'h2a7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2790; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2792 = 10'h2a8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2791; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2793 = 10'h2a9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2792; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2794 = 10'h2aa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2793; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2795 = 10'h2ab == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2794; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2796 = 10'h2ac == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2795; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2797 = 10'h2ad == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2796; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2798 = 10'h2ae == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2797; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2799 = 10'h2af == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2798; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2800 = 10'h2b0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2799; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2801 = 10'h2b1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2800; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2802 = 10'h2b2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2801; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2803 = 10'h2b3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2802; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2804 = 10'h2b4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2803; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2805 = 10'h2b5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2804; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2806 = 10'h2b6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2805; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2807 = 10'h2b7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2806; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2808 = 10'h2b8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2807; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2809 = 10'h2b9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2808; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2810 = 10'h2ba == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2809; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2811 = 10'h2bb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2810; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2812 = 10'h2bc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2811; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2813 = 10'h2bd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2812; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2814 = 10'h2be == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2813; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2815 = 10'h2bf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2814; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2816 = 10'h2c0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2815; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2817 = 10'h2c1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2816; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2818 = 10'h2c2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2817; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2819 = 10'h2c3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2818; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2820 = 10'h2c4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2819; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2821 = 10'h2c5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2820; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2822 = 10'h2c6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2821; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2823 = 10'h2c7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2822; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2824 = 10'h2c8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2823; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2825 = 10'h2c9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2824; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2826 = 10'h2ca == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2825; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2827 = 10'h2cb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2826; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2828 = 10'h2cc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2827; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2829 = 10'h2cd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2828; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2830 = 10'h2ce == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2829; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2831 = 10'h2cf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2830; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2832 = 10'h2d0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2831; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2833 = 10'h2d1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2832; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2834 = 10'h2d2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2833; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2835 = 10'h2d3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2834; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2836 = 10'h2d4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2835; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2837 = 10'h2d5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2836; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2838 = 10'h2d6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2837; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2839 = 10'h2d7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2838; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2840 = 10'h2d8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2839; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2841 = 10'h2d9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2840; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2842 = 10'h2da == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2841; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2843 = 10'h2db == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2842; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2844 = 10'h2dc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2843; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2845 = 10'h2dd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2844; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2846 = 10'h2de == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2845; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2847 = 10'h2df == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2846; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2848 = 10'h2e0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2847; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2849 = 10'h2e1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2848; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2850 = 10'h2e2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2849; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2851 = 10'h2e3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2850; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2852 = 10'h2e4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2851; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2853 = 10'h2e5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2852; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2854 = 10'h2e6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2853; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2855 = 10'h2e7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2854; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2856 = 10'h2e8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2855; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2857 = 10'h2e9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2856; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2858 = 10'h2ea == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2857; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2859 = 10'h2eb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2858; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2860 = 10'h2ec == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2859; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2861 = 10'h2ed == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2860; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2862 = 10'h2ee == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2861; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2863 = 10'h2ef == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2862; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2864 = 10'h2f0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2863; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2865 = 10'h2f1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2864; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2866 = 10'h2f2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2865; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2867 = 10'h2f3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2866; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2868 = 10'h2f4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2867; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2869 = 10'h2f5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2868; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2870 = 10'h2f6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2869; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2871 = 10'h2f7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2870; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2872 = 10'h2f8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2871; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2873 = 10'h2f9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2872; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2874 = 10'h2fa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2873; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2875 = 10'h2fb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2874; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2876 = 10'h2fc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2875; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2877 = 10'h2fd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2876; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2878 = 10'h2fe == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2877; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2879 = 10'h2ff == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2878; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2880 = 10'h300 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2879; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2881 = 10'h301 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2880; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2882 = 10'h302 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2881; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2883 = 10'h303 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2882; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2884 = 10'h304 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2883; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2885 = 10'h305 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2884; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2886 = 10'h306 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2885; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2887 = 10'h307 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2886; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2888 = 10'h308 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2887; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2889 = 10'h309 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2888; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2890 = 10'h30a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2889; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2891 = 10'h30b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2890; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2892 = 10'h30c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2891; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2893 = 10'h30d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2892; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2894 = 10'h30e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2893; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2895 = 10'h30f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2894; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2896 = 10'h310 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2895; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2897 = 10'h311 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2896; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2898 = 10'h312 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2897; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2899 = 10'h313 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2898; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2900 = 10'h314 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2899; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2901 = 10'h315 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2900; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2902 = 10'h316 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2901; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2903 = 10'h317 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2902; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2904 = 10'h318 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2903; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2905 = 10'h319 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2904; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2906 = 10'h31a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2905; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2907 = 10'h31b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2906; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2908 = 10'h31c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2907; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2909 = 10'h31d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2908; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2910 = 10'h31e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2909; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2911 = 10'h31f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2910; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2912 = 10'h320 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2911; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2913 = 10'h321 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2912; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2914 = 10'h322 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2913; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2915 = 10'h323 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2914; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2916 = 10'h324 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2915; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2917 = 10'h325 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2916; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2918 = 10'h326 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2917; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2919 = 10'h327 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2918; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2920 = 10'h328 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2919; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2921 = 10'h329 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2920; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2922 = 10'h32a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2921; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2923 = 10'h32b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2922; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2924 = 10'h32c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2923; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2925 = 10'h32d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2924; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2926 = 10'h32e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2925; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2927 = 10'h32f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2926; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2928 = 10'h330 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2927; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2929 = 10'h331 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2928; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2930 = 10'h332 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2929; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2931 = 10'h333 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2930; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2932 = 10'h334 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2931; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2933 = 10'h335 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2932; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2934 = 10'h336 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2933; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2935 = 10'h337 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2934; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2936 = 10'h338 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2935; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2937 = 10'h339 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2936; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2938 = 10'h33a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2937; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2939 = 10'h33b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2938; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2940 = 10'h33c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2939; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2941 = 10'h33d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2940; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2942 = 10'h33e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2941; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2943 = 10'h33f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2942; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2944 = 10'h340 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2943; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2945 = 10'h341 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2944; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2946 = 10'h342 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2945; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2947 = 10'h343 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2946; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2948 = 10'h344 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2947; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2949 = 10'h345 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2948; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2950 = 10'h346 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2949; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2951 = 10'h347 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2950; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2952 = 10'h348 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2951; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2953 = 10'h349 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2952; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2954 = 10'h34a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2953; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2955 = 10'h34b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2954; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2956 = 10'h34c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2955; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2957 = 10'h34d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2956; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2958 = 10'h34e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2957; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2959 = 10'h34f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2958; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2960 = 10'h350 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2959; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2961 = 10'h351 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2960; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2962 = 10'h352 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2961; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2963 = 10'h353 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2962; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2964 = 10'h354 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2963; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2965 = 10'h355 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2964; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2966 = 10'h356 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2965; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2967 = 10'h357 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2966; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2968 = 10'h358 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2967; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2969 = 10'h359 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2968; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2970 = 10'h35a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2969; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2971 = 10'h35b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2970; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2972 = 10'h35c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2971; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2973 = 10'h35d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2972; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2974 = 10'h35e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2973; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2975 = 10'h35f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2974; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2976 = 10'h360 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2975; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2977 = 10'h361 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2976; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2978 = 10'h362 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2977; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2979 = 10'h363 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2978; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2980 = 10'h364 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2979; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2981 = 10'h365 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2980; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2982 = 10'h366 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2981; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2983 = 10'h367 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2982; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2984 = 10'h368 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2983; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2985 = 10'h369 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2984; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2986 = 10'h36a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2985; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2987 = 10'h36b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2986; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2988 = 10'h36c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2987; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2989 = 10'h36d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2988; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2990 = 10'h36e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2989; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2991 = 10'h36f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2990; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2992 = 10'h370 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2991; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2993 = 10'h371 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2992; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2994 = 10'h372 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2993; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2995 = 10'h373 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2994; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2996 = 10'h374 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2995; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2997 = 10'h375 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2996; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2998 = 10'h376 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2997; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_2999 = 10'h377 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2998; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3000 = 10'h378 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_2999; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3001 = 10'h379 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3000; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3002 = 10'h37a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3001; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3003 = 10'h37b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3002; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3004 = 10'h37c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3003; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3005 = 10'h37d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3004; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3006 = 10'h37e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3005; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3007 = 10'h37f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3006; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3008 = 10'h380 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3007; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3009 = 10'h381 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3008; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3010 = 10'h382 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3009; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3011 = 10'h383 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3010; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3012 = 10'h384 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3011; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3013 = 10'h385 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3012; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3014 = 10'h386 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3013; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3015 = 10'h387 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3014; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3016 = 10'h388 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3015; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3017 = 10'h389 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3016; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3018 = 10'h38a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3017; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3019 = 10'h38b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3018; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3020 = 10'h38c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3019; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3021 = 10'h38d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3020; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3022 = 10'h38e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3021; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3023 = 10'h38f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3022; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3024 = 10'h390 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3023; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3025 = 10'h391 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3024; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3026 = 10'h392 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3025; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3027 = 10'h393 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3026; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3028 = 10'h394 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3027; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3029 = 10'h395 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3028; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3030 = 10'h396 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3029; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3031 = 10'h397 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3030; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3032 = 10'h398 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3031; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3033 = 10'h399 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3032; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3034 = 10'h39a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3033; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3035 = 10'h39b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3034; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3036 = 10'h39c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3035; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3037 = 10'h39d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3036; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3038 = 10'h39e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3037; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3039 = 10'h39f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3038; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3040 = 10'h3a0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3039; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3041 = 10'h3a1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3040; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3042 = 10'h3a2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3041; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3043 = 10'h3a3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3042; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3044 = 10'h3a4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3043; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3045 = 10'h3a5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3044; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3046 = 10'h3a6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3045; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3047 = 10'h3a7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3046; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3048 = 10'h3a8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3047; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3049 = 10'h3a9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3048; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3050 = 10'h3aa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3049; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3051 = 10'h3ab == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3050; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3052 = 10'h3ac == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3051; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3053 = 10'h3ad == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3052; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3054 = 10'h3ae == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3053; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3055 = 10'h3af == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3054; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3056 = 10'h3b0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3055; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3057 = 10'h3b1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3056; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3058 = 10'h3b2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3057; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3059 = 10'h3b3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3058; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3060 = 10'h3b4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3059; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3061 = 10'h3b5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3060; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3062 = 10'h3b6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3061; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3063 = 10'h3b7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3062; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3064 = 10'h3b8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3063; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3065 = 10'h3b9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3064; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3066 = 10'h3ba == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3065; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3067 = 10'h3bb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3066; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3068 = 10'h3bc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3067; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3069 = 10'h3bd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3068; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3070 = 10'h3be == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3069; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3071 = 10'h3bf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3070; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3072 = 10'h3c0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3071; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3073 = 10'h3c1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3072; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3074 = 10'h3c2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3073; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3075 = 10'h3c3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3074; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3076 = 10'h3c4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3075; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3077 = 10'h3c5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3076; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3078 = 10'h3c6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3077; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3079 = 10'h3c7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3078; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3080 = 10'h3c8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3079; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3081 = 10'h3c9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3080; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3082 = 10'h3ca == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3081; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3083 = 10'h3cb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3082; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3084 = 10'h3cc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3083; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3085 = 10'h3cd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3084; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3086 = 10'h3ce == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3085; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3087 = 10'h3cf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3086; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3088 = 10'h3d0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3087; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3089 = 10'h3d1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3088; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3090 = 10'h3d2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3089; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3091 = 10'h3d3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3090; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3092 = 10'h3d4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3091; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3093 = 10'h3d5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3092; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3094 = 10'h3d6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3093; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3095 = 10'h3d7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3094; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3096 = 10'h3d8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3095; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3097 = 10'h3d9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3096; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3098 = 10'h3da == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3097; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3099 = 10'h3db == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3098; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3100 = 10'h3dc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3099; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3101 = 10'h3dd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3100; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3102 = 10'h3de == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3101; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3103 = 10'h3df == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3102; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3104 = 10'h3e0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3103; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3105 = 10'h3e1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3104; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3106 = 10'h3e2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3105; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3107 = 10'h3e3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3106; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3108 = 10'h3e4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3107; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3109 = 10'h3e5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3108; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3110 = 10'h3e6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3109; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3111 = 10'h3e7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3110; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3112 = 10'h3e8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3111; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3113 = 10'h3e9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3112; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3114 = 10'h3ea == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3113; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3115 = 10'h3eb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3114; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3116 = 10'h3ec == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3115; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3117 = 10'h3ed == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3116; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3118 = 10'h3ee == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3117; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3119 = 10'h3ef == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3118; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3120 = 10'h3f0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3119; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3121 = 10'h3f1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3120; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3122 = 10'h3f2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3121; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3123 = 10'h3f3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3122; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3124 = 10'h3f4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3123; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3125 = 10'h3f5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3124; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3126 = 10'h3f6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3125; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3127 = 10'h3f7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3126; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3128 = 10'h3f8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3127; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3129 = 10'h3f9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3128; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3130 = 10'h3fa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3129; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3131 = 10'h3fb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3130; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3132 = 10'h3fc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3131; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3133 = 10'h3fd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3132; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3134 = 10'h3fe == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3133; // @[CPU.scala 125:{16,16}]
  wire [31:0] _GEN_3135 = 10'h3ff == _IFIDIR_T[9:0] ? 32'h0 : _GEN_3134; // @[CPU.scala 125:{16,16}]
  wire [63:0] _PC_T_1 = PC + 64'h4; // @[CPU.scala 126:18]
  wire [12:0] _branchTarget_T_5 = {IFIDIR[31],1'h0,IFIDIR[30:25],IFIDIR[11:7]}; // @[CPU.scala 135:11]
  wire [63:0] _GEN_9496 = {{51{_branchTarget_T_5[12]}},_branchTarget_T_5}; // @[CPU.scala 130:42]
  wire [63:0] branchTarget = $signed(CurPC) + $signed(_GEN_9496); // @[CPU.scala 135:19]
  wire [11:0] _EXMEMALUOut_T_2 = IDEXIR[31:20]; // @[CPU.scala 183:53]
  wire [63:0] _GEN_9497 = {{52{_EXMEMALUOut_T_2[11]}},_EXMEMALUOut_T_2}; // @[CPU.scala 183:36]
  wire [63:0] _EXMEMALUOut_T_6 = $signed(IDEXA) + $signed(_GEN_9497); // @[CPU.scala 183:61]
  wire [11:0] _EXMEMALUOut_T_11 = {IDEXIR[31:25],IDEXrd}; // @[CPU.scala 188:9]
  wire [63:0] _GEN_9498 = {{52{_EXMEMALUOut_T_11[11]}},_EXMEMALUOut_T_11}; // @[CPU.scala 185:36]
  wire [63:0] _EXMEMALUOut_T_15 = $signed(IDEXA) + $signed(_GEN_9498); // @[CPU.scala 188:17]
  wire [31:0] _GEN_3230 = 10'h1 == EXMEMALUOut[9:0] ? DMemory_1 : DMemory_0; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3231 = 10'h2 == EXMEMALUOut[9:0] ? DMemory_2 : _GEN_3230; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3232 = 10'h3 == EXMEMALUOut[9:0] ? DMemory_3 : _GEN_3231; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3233 = 10'h4 == EXMEMALUOut[9:0] ? DMemory_4 : _GEN_3232; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3234 = 10'h5 == EXMEMALUOut[9:0] ? DMemory_5 : _GEN_3233; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3235 = 10'h6 == EXMEMALUOut[9:0] ? DMemory_6 : _GEN_3234; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3236 = 10'h7 == EXMEMALUOut[9:0] ? DMemory_7 : _GEN_3235; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3237 = 10'h8 == EXMEMALUOut[9:0] ? DMemory_8 : _GEN_3236; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3238 = 10'h9 == EXMEMALUOut[9:0] ? DMemory_9 : _GEN_3237; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3239 = 10'ha == EXMEMALUOut[9:0] ? DMemory_10 : _GEN_3238; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3240 = 10'hb == EXMEMALUOut[9:0] ? DMemory_11 : _GEN_3239; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3241 = 10'hc == EXMEMALUOut[9:0] ? DMemory_12 : _GEN_3240; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3242 = 10'hd == EXMEMALUOut[9:0] ? DMemory_13 : _GEN_3241; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3243 = 10'he == EXMEMALUOut[9:0] ? DMemory_14 : _GEN_3242; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3244 = 10'hf == EXMEMALUOut[9:0] ? DMemory_15 : _GEN_3243; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3245 = 10'h10 == EXMEMALUOut[9:0] ? DMemory_16 : _GEN_3244; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3246 = 10'h11 == EXMEMALUOut[9:0] ? DMemory_17 : _GEN_3245; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3247 = 10'h12 == EXMEMALUOut[9:0] ? DMemory_18 : _GEN_3246; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3248 = 10'h13 == EXMEMALUOut[9:0] ? DMemory_19 : _GEN_3247; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3249 = 10'h14 == EXMEMALUOut[9:0] ? DMemory_20 : _GEN_3248; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3250 = 10'h15 == EXMEMALUOut[9:0] ? DMemory_21 : _GEN_3249; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3251 = 10'h16 == EXMEMALUOut[9:0] ? DMemory_22 : _GEN_3250; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3252 = 10'h17 == EXMEMALUOut[9:0] ? DMemory_23 : _GEN_3251; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3253 = 10'h18 == EXMEMALUOut[9:0] ? DMemory_24 : _GEN_3252; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3254 = 10'h19 == EXMEMALUOut[9:0] ? DMemory_25 : _GEN_3253; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3255 = 10'h1a == EXMEMALUOut[9:0] ? DMemory_26 : _GEN_3254; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3256 = 10'h1b == EXMEMALUOut[9:0] ? DMemory_27 : _GEN_3255; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3257 = 10'h1c == EXMEMALUOut[9:0] ? DMemory_28 : _GEN_3256; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3258 = 10'h1d == EXMEMALUOut[9:0] ? DMemory_29 : _GEN_3257; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3259 = 10'h1e == EXMEMALUOut[9:0] ? DMemory_30 : _GEN_3258; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3260 = 10'h1f == EXMEMALUOut[9:0] ? DMemory_31 : _GEN_3259; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3261 = 10'h20 == EXMEMALUOut[9:0] ? DMemory_32 : _GEN_3260; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3262 = 10'h21 == EXMEMALUOut[9:0] ? DMemory_33 : _GEN_3261; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3263 = 10'h22 == EXMEMALUOut[9:0] ? DMemory_34 : _GEN_3262; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3264 = 10'h23 == EXMEMALUOut[9:0] ? DMemory_35 : _GEN_3263; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3265 = 10'h24 == EXMEMALUOut[9:0] ? DMemory_36 : _GEN_3264; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3266 = 10'h25 == EXMEMALUOut[9:0] ? DMemory_37 : _GEN_3265; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3267 = 10'h26 == EXMEMALUOut[9:0] ? DMemory_38 : _GEN_3266; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3268 = 10'h27 == EXMEMALUOut[9:0] ? DMemory_39 : _GEN_3267; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3269 = 10'h28 == EXMEMALUOut[9:0] ? DMemory_40 : _GEN_3268; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3270 = 10'h29 == EXMEMALUOut[9:0] ? DMemory_41 : _GEN_3269; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3271 = 10'h2a == EXMEMALUOut[9:0] ? DMemory_42 : _GEN_3270; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3272 = 10'h2b == EXMEMALUOut[9:0] ? DMemory_43 : _GEN_3271; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3273 = 10'h2c == EXMEMALUOut[9:0] ? DMemory_44 : _GEN_3272; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3274 = 10'h2d == EXMEMALUOut[9:0] ? DMemory_45 : _GEN_3273; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3275 = 10'h2e == EXMEMALUOut[9:0] ? DMemory_46 : _GEN_3274; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3276 = 10'h2f == EXMEMALUOut[9:0] ? DMemory_47 : _GEN_3275; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3277 = 10'h30 == EXMEMALUOut[9:0] ? DMemory_48 : _GEN_3276; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3278 = 10'h31 == EXMEMALUOut[9:0] ? DMemory_49 : _GEN_3277; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3279 = 10'h32 == EXMEMALUOut[9:0] ? DMemory_50 : _GEN_3278; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3280 = 10'h33 == EXMEMALUOut[9:0] ? DMemory_51 : _GEN_3279; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3281 = 10'h34 == EXMEMALUOut[9:0] ? DMemory_52 : _GEN_3280; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3282 = 10'h35 == EXMEMALUOut[9:0] ? DMemory_53 : _GEN_3281; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3283 = 10'h36 == EXMEMALUOut[9:0] ? DMemory_54 : _GEN_3282; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3284 = 10'h37 == EXMEMALUOut[9:0] ? DMemory_55 : _GEN_3283; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3285 = 10'h38 == EXMEMALUOut[9:0] ? DMemory_56 : _GEN_3284; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3286 = 10'h39 == EXMEMALUOut[9:0] ? DMemory_57 : _GEN_3285; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3287 = 10'h3a == EXMEMALUOut[9:0] ? DMemory_58 : _GEN_3286; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3288 = 10'h3b == EXMEMALUOut[9:0] ? DMemory_59 : _GEN_3287; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3289 = 10'h3c == EXMEMALUOut[9:0] ? DMemory_60 : _GEN_3288; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3290 = 10'h3d == EXMEMALUOut[9:0] ? DMemory_61 : _GEN_3289; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3291 = 10'h3e == EXMEMALUOut[9:0] ? DMemory_62 : _GEN_3290; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3292 = 10'h3f == EXMEMALUOut[9:0] ? DMemory_63 : _GEN_3291; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3293 = 10'h40 == EXMEMALUOut[9:0] ? DMemory_64 : _GEN_3292; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3294 = 10'h41 == EXMEMALUOut[9:0] ? DMemory_65 : _GEN_3293; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3295 = 10'h42 == EXMEMALUOut[9:0] ? DMemory_66 : _GEN_3294; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3296 = 10'h43 == EXMEMALUOut[9:0] ? DMemory_67 : _GEN_3295; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3297 = 10'h44 == EXMEMALUOut[9:0] ? DMemory_68 : _GEN_3296; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3298 = 10'h45 == EXMEMALUOut[9:0] ? DMemory_69 : _GEN_3297; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3299 = 10'h46 == EXMEMALUOut[9:0] ? DMemory_70 : _GEN_3298; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3300 = 10'h47 == EXMEMALUOut[9:0] ? DMemory_71 : _GEN_3299; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3301 = 10'h48 == EXMEMALUOut[9:0] ? DMemory_72 : _GEN_3300; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3302 = 10'h49 == EXMEMALUOut[9:0] ? DMemory_73 : _GEN_3301; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3303 = 10'h4a == EXMEMALUOut[9:0] ? DMemory_74 : _GEN_3302; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3304 = 10'h4b == EXMEMALUOut[9:0] ? DMemory_75 : _GEN_3303; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3305 = 10'h4c == EXMEMALUOut[9:0] ? DMemory_76 : _GEN_3304; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3306 = 10'h4d == EXMEMALUOut[9:0] ? DMemory_77 : _GEN_3305; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3307 = 10'h4e == EXMEMALUOut[9:0] ? DMemory_78 : _GEN_3306; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3308 = 10'h4f == EXMEMALUOut[9:0] ? DMemory_79 : _GEN_3307; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3309 = 10'h50 == EXMEMALUOut[9:0] ? DMemory_80 : _GEN_3308; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3310 = 10'h51 == EXMEMALUOut[9:0] ? DMemory_81 : _GEN_3309; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3311 = 10'h52 == EXMEMALUOut[9:0] ? DMemory_82 : _GEN_3310; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3312 = 10'h53 == EXMEMALUOut[9:0] ? DMemory_83 : _GEN_3311; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3313 = 10'h54 == EXMEMALUOut[9:0] ? DMemory_84 : _GEN_3312; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3314 = 10'h55 == EXMEMALUOut[9:0] ? DMemory_85 : _GEN_3313; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3315 = 10'h56 == EXMEMALUOut[9:0] ? DMemory_86 : _GEN_3314; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3316 = 10'h57 == EXMEMALUOut[9:0] ? DMemory_87 : _GEN_3315; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3317 = 10'h58 == EXMEMALUOut[9:0] ? DMemory_88 : _GEN_3316; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3318 = 10'h59 == EXMEMALUOut[9:0] ? DMemory_89 : _GEN_3317; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3319 = 10'h5a == EXMEMALUOut[9:0] ? DMemory_90 : _GEN_3318; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3320 = 10'h5b == EXMEMALUOut[9:0] ? DMemory_91 : _GEN_3319; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3321 = 10'h5c == EXMEMALUOut[9:0] ? DMemory_92 : _GEN_3320; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3322 = 10'h5d == EXMEMALUOut[9:0] ? DMemory_93 : _GEN_3321; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3323 = 10'h5e == EXMEMALUOut[9:0] ? DMemory_94 : _GEN_3322; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3324 = 10'h5f == EXMEMALUOut[9:0] ? DMemory_95 : _GEN_3323; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3325 = 10'h60 == EXMEMALUOut[9:0] ? DMemory_96 : _GEN_3324; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3326 = 10'h61 == EXMEMALUOut[9:0] ? DMemory_97 : _GEN_3325; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3327 = 10'h62 == EXMEMALUOut[9:0] ? DMemory_98 : _GEN_3326; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3328 = 10'h63 == EXMEMALUOut[9:0] ? DMemory_99 : _GEN_3327; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3329 = 10'h64 == EXMEMALUOut[9:0] ? DMemory_100 : _GEN_3328; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3330 = 10'h65 == EXMEMALUOut[9:0] ? DMemory_101 : _GEN_3329; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3331 = 10'h66 == EXMEMALUOut[9:0] ? DMemory_102 : _GEN_3330; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3332 = 10'h67 == EXMEMALUOut[9:0] ? DMemory_103 : _GEN_3331; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3333 = 10'h68 == EXMEMALUOut[9:0] ? DMemory_104 : _GEN_3332; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3334 = 10'h69 == EXMEMALUOut[9:0] ? DMemory_105 : _GEN_3333; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3335 = 10'h6a == EXMEMALUOut[9:0] ? DMemory_106 : _GEN_3334; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3336 = 10'h6b == EXMEMALUOut[9:0] ? DMemory_107 : _GEN_3335; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3337 = 10'h6c == EXMEMALUOut[9:0] ? DMemory_108 : _GEN_3336; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3338 = 10'h6d == EXMEMALUOut[9:0] ? DMemory_109 : _GEN_3337; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3339 = 10'h6e == EXMEMALUOut[9:0] ? DMemory_110 : _GEN_3338; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3340 = 10'h6f == EXMEMALUOut[9:0] ? DMemory_111 : _GEN_3339; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3341 = 10'h70 == EXMEMALUOut[9:0] ? DMemory_112 : _GEN_3340; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3342 = 10'h71 == EXMEMALUOut[9:0] ? DMemory_113 : _GEN_3341; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3343 = 10'h72 == EXMEMALUOut[9:0] ? DMemory_114 : _GEN_3342; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3344 = 10'h73 == EXMEMALUOut[9:0] ? DMemory_115 : _GEN_3343; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3345 = 10'h74 == EXMEMALUOut[9:0] ? DMemory_116 : _GEN_3344; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3346 = 10'h75 == EXMEMALUOut[9:0] ? DMemory_117 : _GEN_3345; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3347 = 10'h76 == EXMEMALUOut[9:0] ? DMemory_118 : _GEN_3346; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3348 = 10'h77 == EXMEMALUOut[9:0] ? DMemory_119 : _GEN_3347; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3349 = 10'h78 == EXMEMALUOut[9:0] ? DMemory_120 : _GEN_3348; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3350 = 10'h79 == EXMEMALUOut[9:0] ? DMemory_121 : _GEN_3349; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3351 = 10'h7a == EXMEMALUOut[9:0] ? DMemory_122 : _GEN_3350; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3352 = 10'h7b == EXMEMALUOut[9:0] ? DMemory_123 : _GEN_3351; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3353 = 10'h7c == EXMEMALUOut[9:0] ? DMemory_124 : _GEN_3352; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3354 = 10'h7d == EXMEMALUOut[9:0] ? DMemory_125 : _GEN_3353; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3355 = 10'h7e == EXMEMALUOut[9:0] ? DMemory_126 : _GEN_3354; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3356 = 10'h7f == EXMEMALUOut[9:0] ? DMemory_127 : _GEN_3355; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3357 = 10'h80 == EXMEMALUOut[9:0] ? DMemory_128 : _GEN_3356; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3358 = 10'h81 == EXMEMALUOut[9:0] ? DMemory_129 : _GEN_3357; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3359 = 10'h82 == EXMEMALUOut[9:0] ? DMemory_130 : _GEN_3358; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3360 = 10'h83 == EXMEMALUOut[9:0] ? DMemory_131 : _GEN_3359; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3361 = 10'h84 == EXMEMALUOut[9:0] ? DMemory_132 : _GEN_3360; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3362 = 10'h85 == EXMEMALUOut[9:0] ? DMemory_133 : _GEN_3361; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3363 = 10'h86 == EXMEMALUOut[9:0] ? DMemory_134 : _GEN_3362; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3364 = 10'h87 == EXMEMALUOut[9:0] ? DMemory_135 : _GEN_3363; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3365 = 10'h88 == EXMEMALUOut[9:0] ? DMemory_136 : _GEN_3364; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3366 = 10'h89 == EXMEMALUOut[9:0] ? DMemory_137 : _GEN_3365; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3367 = 10'h8a == EXMEMALUOut[9:0] ? DMemory_138 : _GEN_3366; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3368 = 10'h8b == EXMEMALUOut[9:0] ? DMemory_139 : _GEN_3367; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3369 = 10'h8c == EXMEMALUOut[9:0] ? DMemory_140 : _GEN_3368; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3370 = 10'h8d == EXMEMALUOut[9:0] ? DMemory_141 : _GEN_3369; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3371 = 10'h8e == EXMEMALUOut[9:0] ? DMemory_142 : _GEN_3370; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3372 = 10'h8f == EXMEMALUOut[9:0] ? DMemory_143 : _GEN_3371; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3373 = 10'h90 == EXMEMALUOut[9:0] ? DMemory_144 : _GEN_3372; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3374 = 10'h91 == EXMEMALUOut[9:0] ? DMemory_145 : _GEN_3373; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3375 = 10'h92 == EXMEMALUOut[9:0] ? DMemory_146 : _GEN_3374; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3376 = 10'h93 == EXMEMALUOut[9:0] ? DMemory_147 : _GEN_3375; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3377 = 10'h94 == EXMEMALUOut[9:0] ? DMemory_148 : _GEN_3376; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3378 = 10'h95 == EXMEMALUOut[9:0] ? DMemory_149 : _GEN_3377; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3379 = 10'h96 == EXMEMALUOut[9:0] ? DMemory_150 : _GEN_3378; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3380 = 10'h97 == EXMEMALUOut[9:0] ? DMemory_151 : _GEN_3379; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3381 = 10'h98 == EXMEMALUOut[9:0] ? DMemory_152 : _GEN_3380; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3382 = 10'h99 == EXMEMALUOut[9:0] ? DMemory_153 : _GEN_3381; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3383 = 10'h9a == EXMEMALUOut[9:0] ? DMemory_154 : _GEN_3382; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3384 = 10'h9b == EXMEMALUOut[9:0] ? DMemory_155 : _GEN_3383; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3385 = 10'h9c == EXMEMALUOut[9:0] ? DMemory_156 : _GEN_3384; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3386 = 10'h9d == EXMEMALUOut[9:0] ? DMemory_157 : _GEN_3385; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3387 = 10'h9e == EXMEMALUOut[9:0] ? DMemory_158 : _GEN_3386; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3388 = 10'h9f == EXMEMALUOut[9:0] ? DMemory_159 : _GEN_3387; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3389 = 10'ha0 == EXMEMALUOut[9:0] ? DMemory_160 : _GEN_3388; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3390 = 10'ha1 == EXMEMALUOut[9:0] ? DMemory_161 : _GEN_3389; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3391 = 10'ha2 == EXMEMALUOut[9:0] ? DMemory_162 : _GEN_3390; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3392 = 10'ha3 == EXMEMALUOut[9:0] ? DMemory_163 : _GEN_3391; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3393 = 10'ha4 == EXMEMALUOut[9:0] ? DMemory_164 : _GEN_3392; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3394 = 10'ha5 == EXMEMALUOut[9:0] ? DMemory_165 : _GEN_3393; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3395 = 10'ha6 == EXMEMALUOut[9:0] ? DMemory_166 : _GEN_3394; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3396 = 10'ha7 == EXMEMALUOut[9:0] ? DMemory_167 : _GEN_3395; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3397 = 10'ha8 == EXMEMALUOut[9:0] ? DMemory_168 : _GEN_3396; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3398 = 10'ha9 == EXMEMALUOut[9:0] ? DMemory_169 : _GEN_3397; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3399 = 10'haa == EXMEMALUOut[9:0] ? DMemory_170 : _GEN_3398; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3400 = 10'hab == EXMEMALUOut[9:0] ? DMemory_171 : _GEN_3399; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3401 = 10'hac == EXMEMALUOut[9:0] ? DMemory_172 : _GEN_3400; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3402 = 10'had == EXMEMALUOut[9:0] ? DMemory_173 : _GEN_3401; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3403 = 10'hae == EXMEMALUOut[9:0] ? DMemory_174 : _GEN_3402; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3404 = 10'haf == EXMEMALUOut[9:0] ? DMemory_175 : _GEN_3403; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3405 = 10'hb0 == EXMEMALUOut[9:0] ? DMemory_176 : _GEN_3404; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3406 = 10'hb1 == EXMEMALUOut[9:0] ? DMemory_177 : _GEN_3405; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3407 = 10'hb2 == EXMEMALUOut[9:0] ? DMemory_178 : _GEN_3406; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3408 = 10'hb3 == EXMEMALUOut[9:0] ? DMemory_179 : _GEN_3407; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3409 = 10'hb4 == EXMEMALUOut[9:0] ? DMemory_180 : _GEN_3408; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3410 = 10'hb5 == EXMEMALUOut[9:0] ? DMemory_181 : _GEN_3409; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3411 = 10'hb6 == EXMEMALUOut[9:0] ? DMemory_182 : _GEN_3410; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3412 = 10'hb7 == EXMEMALUOut[9:0] ? DMemory_183 : _GEN_3411; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3413 = 10'hb8 == EXMEMALUOut[9:0] ? DMemory_184 : _GEN_3412; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3414 = 10'hb9 == EXMEMALUOut[9:0] ? DMemory_185 : _GEN_3413; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3415 = 10'hba == EXMEMALUOut[9:0] ? DMemory_186 : _GEN_3414; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3416 = 10'hbb == EXMEMALUOut[9:0] ? DMemory_187 : _GEN_3415; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3417 = 10'hbc == EXMEMALUOut[9:0] ? DMemory_188 : _GEN_3416; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3418 = 10'hbd == EXMEMALUOut[9:0] ? DMemory_189 : _GEN_3417; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3419 = 10'hbe == EXMEMALUOut[9:0] ? DMemory_190 : _GEN_3418; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3420 = 10'hbf == EXMEMALUOut[9:0] ? DMemory_191 : _GEN_3419; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3421 = 10'hc0 == EXMEMALUOut[9:0] ? DMemory_192 : _GEN_3420; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3422 = 10'hc1 == EXMEMALUOut[9:0] ? DMemory_193 : _GEN_3421; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3423 = 10'hc2 == EXMEMALUOut[9:0] ? DMemory_194 : _GEN_3422; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3424 = 10'hc3 == EXMEMALUOut[9:0] ? DMemory_195 : _GEN_3423; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3425 = 10'hc4 == EXMEMALUOut[9:0] ? DMemory_196 : _GEN_3424; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3426 = 10'hc5 == EXMEMALUOut[9:0] ? DMemory_197 : _GEN_3425; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3427 = 10'hc6 == EXMEMALUOut[9:0] ? DMemory_198 : _GEN_3426; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3428 = 10'hc7 == EXMEMALUOut[9:0] ? DMemory_199 : _GEN_3427; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3429 = 10'hc8 == EXMEMALUOut[9:0] ? DMemory_200 : _GEN_3428; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3430 = 10'hc9 == EXMEMALUOut[9:0] ? DMemory_201 : _GEN_3429; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3431 = 10'hca == EXMEMALUOut[9:0] ? DMemory_202 : _GEN_3430; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3432 = 10'hcb == EXMEMALUOut[9:0] ? DMemory_203 : _GEN_3431; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3433 = 10'hcc == EXMEMALUOut[9:0] ? DMemory_204 : _GEN_3432; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3434 = 10'hcd == EXMEMALUOut[9:0] ? DMemory_205 : _GEN_3433; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3435 = 10'hce == EXMEMALUOut[9:0] ? DMemory_206 : _GEN_3434; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3436 = 10'hcf == EXMEMALUOut[9:0] ? DMemory_207 : _GEN_3435; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3437 = 10'hd0 == EXMEMALUOut[9:0] ? DMemory_208 : _GEN_3436; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3438 = 10'hd1 == EXMEMALUOut[9:0] ? DMemory_209 : _GEN_3437; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3439 = 10'hd2 == EXMEMALUOut[9:0] ? DMemory_210 : _GEN_3438; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3440 = 10'hd3 == EXMEMALUOut[9:0] ? DMemory_211 : _GEN_3439; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3441 = 10'hd4 == EXMEMALUOut[9:0] ? DMemory_212 : _GEN_3440; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3442 = 10'hd5 == EXMEMALUOut[9:0] ? DMemory_213 : _GEN_3441; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3443 = 10'hd6 == EXMEMALUOut[9:0] ? DMemory_214 : _GEN_3442; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3444 = 10'hd7 == EXMEMALUOut[9:0] ? DMemory_215 : _GEN_3443; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3445 = 10'hd8 == EXMEMALUOut[9:0] ? DMemory_216 : _GEN_3444; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3446 = 10'hd9 == EXMEMALUOut[9:0] ? DMemory_217 : _GEN_3445; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3447 = 10'hda == EXMEMALUOut[9:0] ? DMemory_218 : _GEN_3446; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3448 = 10'hdb == EXMEMALUOut[9:0] ? DMemory_219 : _GEN_3447; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3449 = 10'hdc == EXMEMALUOut[9:0] ? DMemory_220 : _GEN_3448; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3450 = 10'hdd == EXMEMALUOut[9:0] ? DMemory_221 : _GEN_3449; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3451 = 10'hde == EXMEMALUOut[9:0] ? DMemory_222 : _GEN_3450; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3452 = 10'hdf == EXMEMALUOut[9:0] ? DMemory_223 : _GEN_3451; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3453 = 10'he0 == EXMEMALUOut[9:0] ? DMemory_224 : _GEN_3452; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3454 = 10'he1 == EXMEMALUOut[9:0] ? DMemory_225 : _GEN_3453; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3455 = 10'he2 == EXMEMALUOut[9:0] ? DMemory_226 : _GEN_3454; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3456 = 10'he3 == EXMEMALUOut[9:0] ? DMemory_227 : _GEN_3455; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3457 = 10'he4 == EXMEMALUOut[9:0] ? DMemory_228 : _GEN_3456; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3458 = 10'he5 == EXMEMALUOut[9:0] ? DMemory_229 : _GEN_3457; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3459 = 10'he6 == EXMEMALUOut[9:0] ? DMemory_230 : _GEN_3458; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3460 = 10'he7 == EXMEMALUOut[9:0] ? DMemory_231 : _GEN_3459; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3461 = 10'he8 == EXMEMALUOut[9:0] ? DMemory_232 : _GEN_3460; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3462 = 10'he9 == EXMEMALUOut[9:0] ? DMemory_233 : _GEN_3461; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3463 = 10'hea == EXMEMALUOut[9:0] ? DMemory_234 : _GEN_3462; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3464 = 10'heb == EXMEMALUOut[9:0] ? DMemory_235 : _GEN_3463; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3465 = 10'hec == EXMEMALUOut[9:0] ? DMemory_236 : _GEN_3464; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3466 = 10'hed == EXMEMALUOut[9:0] ? DMemory_237 : _GEN_3465; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3467 = 10'hee == EXMEMALUOut[9:0] ? DMemory_238 : _GEN_3466; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3468 = 10'hef == EXMEMALUOut[9:0] ? DMemory_239 : _GEN_3467; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3469 = 10'hf0 == EXMEMALUOut[9:0] ? DMemory_240 : _GEN_3468; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3470 = 10'hf1 == EXMEMALUOut[9:0] ? DMemory_241 : _GEN_3469; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3471 = 10'hf2 == EXMEMALUOut[9:0] ? DMemory_242 : _GEN_3470; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3472 = 10'hf3 == EXMEMALUOut[9:0] ? DMemory_243 : _GEN_3471; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3473 = 10'hf4 == EXMEMALUOut[9:0] ? DMemory_244 : _GEN_3472; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3474 = 10'hf5 == EXMEMALUOut[9:0] ? DMemory_245 : _GEN_3473; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3475 = 10'hf6 == EXMEMALUOut[9:0] ? DMemory_246 : _GEN_3474; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3476 = 10'hf7 == EXMEMALUOut[9:0] ? DMemory_247 : _GEN_3475; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3477 = 10'hf8 == EXMEMALUOut[9:0] ? DMemory_248 : _GEN_3476; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3478 = 10'hf9 == EXMEMALUOut[9:0] ? DMemory_249 : _GEN_3477; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3479 = 10'hfa == EXMEMALUOut[9:0] ? DMemory_250 : _GEN_3478; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3480 = 10'hfb == EXMEMALUOut[9:0] ? DMemory_251 : _GEN_3479; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3481 = 10'hfc == EXMEMALUOut[9:0] ? DMemory_252 : _GEN_3480; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3482 = 10'hfd == EXMEMALUOut[9:0] ? DMemory_253 : _GEN_3481; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3483 = 10'hfe == EXMEMALUOut[9:0] ? DMemory_254 : _GEN_3482; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3484 = 10'hff == EXMEMALUOut[9:0] ? DMemory_255 : _GEN_3483; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3485 = 10'h100 == EXMEMALUOut[9:0] ? DMemory_256 : _GEN_3484; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3486 = 10'h101 == EXMEMALUOut[9:0] ? DMemory_257 : _GEN_3485; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3487 = 10'h102 == EXMEMALUOut[9:0] ? DMemory_258 : _GEN_3486; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3488 = 10'h103 == EXMEMALUOut[9:0] ? DMemory_259 : _GEN_3487; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3489 = 10'h104 == EXMEMALUOut[9:0] ? DMemory_260 : _GEN_3488; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3490 = 10'h105 == EXMEMALUOut[9:0] ? DMemory_261 : _GEN_3489; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3491 = 10'h106 == EXMEMALUOut[9:0] ? DMemory_262 : _GEN_3490; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3492 = 10'h107 == EXMEMALUOut[9:0] ? DMemory_263 : _GEN_3491; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3493 = 10'h108 == EXMEMALUOut[9:0] ? DMemory_264 : _GEN_3492; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3494 = 10'h109 == EXMEMALUOut[9:0] ? DMemory_265 : _GEN_3493; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3495 = 10'h10a == EXMEMALUOut[9:0] ? DMemory_266 : _GEN_3494; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3496 = 10'h10b == EXMEMALUOut[9:0] ? DMemory_267 : _GEN_3495; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3497 = 10'h10c == EXMEMALUOut[9:0] ? DMemory_268 : _GEN_3496; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3498 = 10'h10d == EXMEMALUOut[9:0] ? DMemory_269 : _GEN_3497; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3499 = 10'h10e == EXMEMALUOut[9:0] ? DMemory_270 : _GEN_3498; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3500 = 10'h10f == EXMEMALUOut[9:0] ? DMemory_271 : _GEN_3499; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3501 = 10'h110 == EXMEMALUOut[9:0] ? DMemory_272 : _GEN_3500; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3502 = 10'h111 == EXMEMALUOut[9:0] ? DMemory_273 : _GEN_3501; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3503 = 10'h112 == EXMEMALUOut[9:0] ? DMemory_274 : _GEN_3502; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3504 = 10'h113 == EXMEMALUOut[9:0] ? DMemory_275 : _GEN_3503; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3505 = 10'h114 == EXMEMALUOut[9:0] ? DMemory_276 : _GEN_3504; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3506 = 10'h115 == EXMEMALUOut[9:0] ? DMemory_277 : _GEN_3505; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3507 = 10'h116 == EXMEMALUOut[9:0] ? DMemory_278 : _GEN_3506; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3508 = 10'h117 == EXMEMALUOut[9:0] ? DMemory_279 : _GEN_3507; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3509 = 10'h118 == EXMEMALUOut[9:0] ? DMemory_280 : _GEN_3508; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3510 = 10'h119 == EXMEMALUOut[9:0] ? DMemory_281 : _GEN_3509; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3511 = 10'h11a == EXMEMALUOut[9:0] ? DMemory_282 : _GEN_3510; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3512 = 10'h11b == EXMEMALUOut[9:0] ? DMemory_283 : _GEN_3511; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3513 = 10'h11c == EXMEMALUOut[9:0] ? DMemory_284 : _GEN_3512; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3514 = 10'h11d == EXMEMALUOut[9:0] ? DMemory_285 : _GEN_3513; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3515 = 10'h11e == EXMEMALUOut[9:0] ? DMemory_286 : _GEN_3514; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3516 = 10'h11f == EXMEMALUOut[9:0] ? DMemory_287 : _GEN_3515; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3517 = 10'h120 == EXMEMALUOut[9:0] ? DMemory_288 : _GEN_3516; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3518 = 10'h121 == EXMEMALUOut[9:0] ? DMemory_289 : _GEN_3517; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3519 = 10'h122 == EXMEMALUOut[9:0] ? DMemory_290 : _GEN_3518; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3520 = 10'h123 == EXMEMALUOut[9:0] ? DMemory_291 : _GEN_3519; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3521 = 10'h124 == EXMEMALUOut[9:0] ? DMemory_292 : _GEN_3520; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3522 = 10'h125 == EXMEMALUOut[9:0] ? DMemory_293 : _GEN_3521; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3523 = 10'h126 == EXMEMALUOut[9:0] ? DMemory_294 : _GEN_3522; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3524 = 10'h127 == EXMEMALUOut[9:0] ? DMemory_295 : _GEN_3523; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3525 = 10'h128 == EXMEMALUOut[9:0] ? DMemory_296 : _GEN_3524; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3526 = 10'h129 == EXMEMALUOut[9:0] ? DMemory_297 : _GEN_3525; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3527 = 10'h12a == EXMEMALUOut[9:0] ? DMemory_298 : _GEN_3526; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3528 = 10'h12b == EXMEMALUOut[9:0] ? DMemory_299 : _GEN_3527; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3529 = 10'h12c == EXMEMALUOut[9:0] ? DMemory_300 : _GEN_3528; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3530 = 10'h12d == EXMEMALUOut[9:0] ? DMemory_301 : _GEN_3529; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3531 = 10'h12e == EXMEMALUOut[9:0] ? DMemory_302 : _GEN_3530; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3532 = 10'h12f == EXMEMALUOut[9:0] ? DMemory_303 : _GEN_3531; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3533 = 10'h130 == EXMEMALUOut[9:0] ? DMemory_304 : _GEN_3532; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3534 = 10'h131 == EXMEMALUOut[9:0] ? DMemory_305 : _GEN_3533; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3535 = 10'h132 == EXMEMALUOut[9:0] ? DMemory_306 : _GEN_3534; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3536 = 10'h133 == EXMEMALUOut[9:0] ? DMemory_307 : _GEN_3535; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3537 = 10'h134 == EXMEMALUOut[9:0] ? DMemory_308 : _GEN_3536; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3538 = 10'h135 == EXMEMALUOut[9:0] ? DMemory_309 : _GEN_3537; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3539 = 10'h136 == EXMEMALUOut[9:0] ? DMemory_310 : _GEN_3538; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3540 = 10'h137 == EXMEMALUOut[9:0] ? DMemory_311 : _GEN_3539; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3541 = 10'h138 == EXMEMALUOut[9:0] ? DMemory_312 : _GEN_3540; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3542 = 10'h139 == EXMEMALUOut[9:0] ? DMemory_313 : _GEN_3541; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3543 = 10'h13a == EXMEMALUOut[9:0] ? DMemory_314 : _GEN_3542; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3544 = 10'h13b == EXMEMALUOut[9:0] ? DMemory_315 : _GEN_3543; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3545 = 10'h13c == EXMEMALUOut[9:0] ? DMemory_316 : _GEN_3544; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3546 = 10'h13d == EXMEMALUOut[9:0] ? DMemory_317 : _GEN_3545; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3547 = 10'h13e == EXMEMALUOut[9:0] ? DMemory_318 : _GEN_3546; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3548 = 10'h13f == EXMEMALUOut[9:0] ? DMemory_319 : _GEN_3547; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3549 = 10'h140 == EXMEMALUOut[9:0] ? DMemory_320 : _GEN_3548; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3550 = 10'h141 == EXMEMALUOut[9:0] ? DMemory_321 : _GEN_3549; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3551 = 10'h142 == EXMEMALUOut[9:0] ? DMemory_322 : _GEN_3550; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3552 = 10'h143 == EXMEMALUOut[9:0] ? DMemory_323 : _GEN_3551; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3553 = 10'h144 == EXMEMALUOut[9:0] ? DMemory_324 : _GEN_3552; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3554 = 10'h145 == EXMEMALUOut[9:0] ? DMemory_325 : _GEN_3553; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3555 = 10'h146 == EXMEMALUOut[9:0] ? DMemory_326 : _GEN_3554; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3556 = 10'h147 == EXMEMALUOut[9:0] ? DMemory_327 : _GEN_3555; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3557 = 10'h148 == EXMEMALUOut[9:0] ? DMemory_328 : _GEN_3556; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3558 = 10'h149 == EXMEMALUOut[9:0] ? DMemory_329 : _GEN_3557; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3559 = 10'h14a == EXMEMALUOut[9:0] ? DMemory_330 : _GEN_3558; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3560 = 10'h14b == EXMEMALUOut[9:0] ? DMemory_331 : _GEN_3559; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3561 = 10'h14c == EXMEMALUOut[9:0] ? DMemory_332 : _GEN_3560; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3562 = 10'h14d == EXMEMALUOut[9:0] ? DMemory_333 : _GEN_3561; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3563 = 10'h14e == EXMEMALUOut[9:0] ? DMemory_334 : _GEN_3562; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3564 = 10'h14f == EXMEMALUOut[9:0] ? DMemory_335 : _GEN_3563; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3565 = 10'h150 == EXMEMALUOut[9:0] ? DMemory_336 : _GEN_3564; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3566 = 10'h151 == EXMEMALUOut[9:0] ? DMemory_337 : _GEN_3565; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3567 = 10'h152 == EXMEMALUOut[9:0] ? DMemory_338 : _GEN_3566; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3568 = 10'h153 == EXMEMALUOut[9:0] ? DMemory_339 : _GEN_3567; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3569 = 10'h154 == EXMEMALUOut[9:0] ? DMemory_340 : _GEN_3568; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3570 = 10'h155 == EXMEMALUOut[9:0] ? DMemory_341 : _GEN_3569; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3571 = 10'h156 == EXMEMALUOut[9:0] ? DMemory_342 : _GEN_3570; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3572 = 10'h157 == EXMEMALUOut[9:0] ? DMemory_343 : _GEN_3571; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3573 = 10'h158 == EXMEMALUOut[9:0] ? DMemory_344 : _GEN_3572; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3574 = 10'h159 == EXMEMALUOut[9:0] ? DMemory_345 : _GEN_3573; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3575 = 10'h15a == EXMEMALUOut[9:0] ? DMemory_346 : _GEN_3574; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3576 = 10'h15b == EXMEMALUOut[9:0] ? DMemory_347 : _GEN_3575; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3577 = 10'h15c == EXMEMALUOut[9:0] ? DMemory_348 : _GEN_3576; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3578 = 10'h15d == EXMEMALUOut[9:0] ? DMemory_349 : _GEN_3577; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3579 = 10'h15e == EXMEMALUOut[9:0] ? DMemory_350 : _GEN_3578; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3580 = 10'h15f == EXMEMALUOut[9:0] ? DMemory_351 : _GEN_3579; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3581 = 10'h160 == EXMEMALUOut[9:0] ? DMemory_352 : _GEN_3580; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3582 = 10'h161 == EXMEMALUOut[9:0] ? DMemory_353 : _GEN_3581; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3583 = 10'h162 == EXMEMALUOut[9:0] ? DMemory_354 : _GEN_3582; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3584 = 10'h163 == EXMEMALUOut[9:0] ? DMemory_355 : _GEN_3583; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3585 = 10'h164 == EXMEMALUOut[9:0] ? DMemory_356 : _GEN_3584; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3586 = 10'h165 == EXMEMALUOut[9:0] ? DMemory_357 : _GEN_3585; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3587 = 10'h166 == EXMEMALUOut[9:0] ? DMemory_358 : _GEN_3586; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3588 = 10'h167 == EXMEMALUOut[9:0] ? DMemory_359 : _GEN_3587; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3589 = 10'h168 == EXMEMALUOut[9:0] ? DMemory_360 : _GEN_3588; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3590 = 10'h169 == EXMEMALUOut[9:0] ? DMemory_361 : _GEN_3589; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3591 = 10'h16a == EXMEMALUOut[9:0] ? DMemory_362 : _GEN_3590; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3592 = 10'h16b == EXMEMALUOut[9:0] ? DMemory_363 : _GEN_3591; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3593 = 10'h16c == EXMEMALUOut[9:0] ? DMemory_364 : _GEN_3592; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3594 = 10'h16d == EXMEMALUOut[9:0] ? DMemory_365 : _GEN_3593; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3595 = 10'h16e == EXMEMALUOut[9:0] ? DMemory_366 : _GEN_3594; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3596 = 10'h16f == EXMEMALUOut[9:0] ? DMemory_367 : _GEN_3595; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3597 = 10'h170 == EXMEMALUOut[9:0] ? DMemory_368 : _GEN_3596; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3598 = 10'h171 == EXMEMALUOut[9:0] ? DMemory_369 : _GEN_3597; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3599 = 10'h172 == EXMEMALUOut[9:0] ? DMemory_370 : _GEN_3598; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3600 = 10'h173 == EXMEMALUOut[9:0] ? DMemory_371 : _GEN_3599; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3601 = 10'h174 == EXMEMALUOut[9:0] ? DMemory_372 : _GEN_3600; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3602 = 10'h175 == EXMEMALUOut[9:0] ? DMemory_373 : _GEN_3601; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3603 = 10'h176 == EXMEMALUOut[9:0] ? DMemory_374 : _GEN_3602; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3604 = 10'h177 == EXMEMALUOut[9:0] ? DMemory_375 : _GEN_3603; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3605 = 10'h178 == EXMEMALUOut[9:0] ? DMemory_376 : _GEN_3604; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3606 = 10'h179 == EXMEMALUOut[9:0] ? DMemory_377 : _GEN_3605; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3607 = 10'h17a == EXMEMALUOut[9:0] ? DMemory_378 : _GEN_3606; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3608 = 10'h17b == EXMEMALUOut[9:0] ? DMemory_379 : _GEN_3607; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3609 = 10'h17c == EXMEMALUOut[9:0] ? DMemory_380 : _GEN_3608; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3610 = 10'h17d == EXMEMALUOut[9:0] ? DMemory_381 : _GEN_3609; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3611 = 10'h17e == EXMEMALUOut[9:0] ? DMemory_382 : _GEN_3610; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3612 = 10'h17f == EXMEMALUOut[9:0] ? DMemory_383 : _GEN_3611; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3613 = 10'h180 == EXMEMALUOut[9:0] ? DMemory_384 : _GEN_3612; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3614 = 10'h181 == EXMEMALUOut[9:0] ? DMemory_385 : _GEN_3613; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3615 = 10'h182 == EXMEMALUOut[9:0] ? DMemory_386 : _GEN_3614; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3616 = 10'h183 == EXMEMALUOut[9:0] ? DMemory_387 : _GEN_3615; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3617 = 10'h184 == EXMEMALUOut[9:0] ? DMemory_388 : _GEN_3616; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3618 = 10'h185 == EXMEMALUOut[9:0] ? DMemory_389 : _GEN_3617; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3619 = 10'h186 == EXMEMALUOut[9:0] ? DMemory_390 : _GEN_3618; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3620 = 10'h187 == EXMEMALUOut[9:0] ? DMemory_391 : _GEN_3619; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3621 = 10'h188 == EXMEMALUOut[9:0] ? DMemory_392 : _GEN_3620; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3622 = 10'h189 == EXMEMALUOut[9:0] ? DMemory_393 : _GEN_3621; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3623 = 10'h18a == EXMEMALUOut[9:0] ? DMemory_394 : _GEN_3622; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3624 = 10'h18b == EXMEMALUOut[9:0] ? DMemory_395 : _GEN_3623; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3625 = 10'h18c == EXMEMALUOut[9:0] ? DMemory_396 : _GEN_3624; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3626 = 10'h18d == EXMEMALUOut[9:0] ? DMemory_397 : _GEN_3625; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3627 = 10'h18e == EXMEMALUOut[9:0] ? DMemory_398 : _GEN_3626; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3628 = 10'h18f == EXMEMALUOut[9:0] ? DMemory_399 : _GEN_3627; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3629 = 10'h190 == EXMEMALUOut[9:0] ? DMemory_400 : _GEN_3628; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3630 = 10'h191 == EXMEMALUOut[9:0] ? DMemory_401 : _GEN_3629; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3631 = 10'h192 == EXMEMALUOut[9:0] ? DMemory_402 : _GEN_3630; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3632 = 10'h193 == EXMEMALUOut[9:0] ? DMemory_403 : _GEN_3631; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3633 = 10'h194 == EXMEMALUOut[9:0] ? DMemory_404 : _GEN_3632; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3634 = 10'h195 == EXMEMALUOut[9:0] ? DMemory_405 : _GEN_3633; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3635 = 10'h196 == EXMEMALUOut[9:0] ? DMemory_406 : _GEN_3634; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3636 = 10'h197 == EXMEMALUOut[9:0] ? DMemory_407 : _GEN_3635; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3637 = 10'h198 == EXMEMALUOut[9:0] ? DMemory_408 : _GEN_3636; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3638 = 10'h199 == EXMEMALUOut[9:0] ? DMemory_409 : _GEN_3637; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3639 = 10'h19a == EXMEMALUOut[9:0] ? DMemory_410 : _GEN_3638; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3640 = 10'h19b == EXMEMALUOut[9:0] ? DMemory_411 : _GEN_3639; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3641 = 10'h19c == EXMEMALUOut[9:0] ? DMemory_412 : _GEN_3640; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3642 = 10'h19d == EXMEMALUOut[9:0] ? DMemory_413 : _GEN_3641; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3643 = 10'h19e == EXMEMALUOut[9:0] ? DMemory_414 : _GEN_3642; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3644 = 10'h19f == EXMEMALUOut[9:0] ? DMemory_415 : _GEN_3643; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3645 = 10'h1a0 == EXMEMALUOut[9:0] ? DMemory_416 : _GEN_3644; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3646 = 10'h1a1 == EXMEMALUOut[9:0] ? DMemory_417 : _GEN_3645; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3647 = 10'h1a2 == EXMEMALUOut[9:0] ? DMemory_418 : _GEN_3646; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3648 = 10'h1a3 == EXMEMALUOut[9:0] ? DMemory_419 : _GEN_3647; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3649 = 10'h1a4 == EXMEMALUOut[9:0] ? DMemory_420 : _GEN_3648; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3650 = 10'h1a5 == EXMEMALUOut[9:0] ? DMemory_421 : _GEN_3649; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3651 = 10'h1a6 == EXMEMALUOut[9:0] ? DMemory_422 : _GEN_3650; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3652 = 10'h1a7 == EXMEMALUOut[9:0] ? DMemory_423 : _GEN_3651; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3653 = 10'h1a8 == EXMEMALUOut[9:0] ? DMemory_424 : _GEN_3652; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3654 = 10'h1a9 == EXMEMALUOut[9:0] ? DMemory_425 : _GEN_3653; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3655 = 10'h1aa == EXMEMALUOut[9:0] ? DMemory_426 : _GEN_3654; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3656 = 10'h1ab == EXMEMALUOut[9:0] ? DMemory_427 : _GEN_3655; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3657 = 10'h1ac == EXMEMALUOut[9:0] ? DMemory_428 : _GEN_3656; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3658 = 10'h1ad == EXMEMALUOut[9:0] ? DMemory_429 : _GEN_3657; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3659 = 10'h1ae == EXMEMALUOut[9:0] ? DMemory_430 : _GEN_3658; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3660 = 10'h1af == EXMEMALUOut[9:0] ? DMemory_431 : _GEN_3659; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3661 = 10'h1b0 == EXMEMALUOut[9:0] ? DMemory_432 : _GEN_3660; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3662 = 10'h1b1 == EXMEMALUOut[9:0] ? DMemory_433 : _GEN_3661; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3663 = 10'h1b2 == EXMEMALUOut[9:0] ? DMemory_434 : _GEN_3662; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3664 = 10'h1b3 == EXMEMALUOut[9:0] ? DMemory_435 : _GEN_3663; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3665 = 10'h1b4 == EXMEMALUOut[9:0] ? DMemory_436 : _GEN_3664; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3666 = 10'h1b5 == EXMEMALUOut[9:0] ? DMemory_437 : _GEN_3665; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3667 = 10'h1b6 == EXMEMALUOut[9:0] ? DMemory_438 : _GEN_3666; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3668 = 10'h1b7 == EXMEMALUOut[9:0] ? DMemory_439 : _GEN_3667; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3669 = 10'h1b8 == EXMEMALUOut[9:0] ? DMemory_440 : _GEN_3668; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3670 = 10'h1b9 == EXMEMALUOut[9:0] ? DMemory_441 : _GEN_3669; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3671 = 10'h1ba == EXMEMALUOut[9:0] ? DMemory_442 : _GEN_3670; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3672 = 10'h1bb == EXMEMALUOut[9:0] ? DMemory_443 : _GEN_3671; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3673 = 10'h1bc == EXMEMALUOut[9:0] ? DMemory_444 : _GEN_3672; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3674 = 10'h1bd == EXMEMALUOut[9:0] ? DMemory_445 : _GEN_3673; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3675 = 10'h1be == EXMEMALUOut[9:0] ? DMemory_446 : _GEN_3674; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3676 = 10'h1bf == EXMEMALUOut[9:0] ? DMemory_447 : _GEN_3675; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3677 = 10'h1c0 == EXMEMALUOut[9:0] ? DMemory_448 : _GEN_3676; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3678 = 10'h1c1 == EXMEMALUOut[9:0] ? DMemory_449 : _GEN_3677; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3679 = 10'h1c2 == EXMEMALUOut[9:0] ? DMemory_450 : _GEN_3678; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3680 = 10'h1c3 == EXMEMALUOut[9:0] ? DMemory_451 : _GEN_3679; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3681 = 10'h1c4 == EXMEMALUOut[9:0] ? DMemory_452 : _GEN_3680; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3682 = 10'h1c5 == EXMEMALUOut[9:0] ? DMemory_453 : _GEN_3681; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3683 = 10'h1c6 == EXMEMALUOut[9:0] ? DMemory_454 : _GEN_3682; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3684 = 10'h1c7 == EXMEMALUOut[9:0] ? DMemory_455 : _GEN_3683; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3685 = 10'h1c8 == EXMEMALUOut[9:0] ? DMemory_456 : _GEN_3684; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3686 = 10'h1c9 == EXMEMALUOut[9:0] ? DMemory_457 : _GEN_3685; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3687 = 10'h1ca == EXMEMALUOut[9:0] ? DMemory_458 : _GEN_3686; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3688 = 10'h1cb == EXMEMALUOut[9:0] ? DMemory_459 : _GEN_3687; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3689 = 10'h1cc == EXMEMALUOut[9:0] ? DMemory_460 : _GEN_3688; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3690 = 10'h1cd == EXMEMALUOut[9:0] ? DMemory_461 : _GEN_3689; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3691 = 10'h1ce == EXMEMALUOut[9:0] ? DMemory_462 : _GEN_3690; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3692 = 10'h1cf == EXMEMALUOut[9:0] ? DMemory_463 : _GEN_3691; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3693 = 10'h1d0 == EXMEMALUOut[9:0] ? DMemory_464 : _GEN_3692; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3694 = 10'h1d1 == EXMEMALUOut[9:0] ? DMemory_465 : _GEN_3693; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3695 = 10'h1d2 == EXMEMALUOut[9:0] ? DMemory_466 : _GEN_3694; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3696 = 10'h1d3 == EXMEMALUOut[9:0] ? DMemory_467 : _GEN_3695; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3697 = 10'h1d4 == EXMEMALUOut[9:0] ? DMemory_468 : _GEN_3696; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3698 = 10'h1d5 == EXMEMALUOut[9:0] ? DMemory_469 : _GEN_3697; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3699 = 10'h1d6 == EXMEMALUOut[9:0] ? DMemory_470 : _GEN_3698; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3700 = 10'h1d7 == EXMEMALUOut[9:0] ? DMemory_471 : _GEN_3699; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3701 = 10'h1d8 == EXMEMALUOut[9:0] ? DMemory_472 : _GEN_3700; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3702 = 10'h1d9 == EXMEMALUOut[9:0] ? DMemory_473 : _GEN_3701; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3703 = 10'h1da == EXMEMALUOut[9:0] ? DMemory_474 : _GEN_3702; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3704 = 10'h1db == EXMEMALUOut[9:0] ? DMemory_475 : _GEN_3703; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3705 = 10'h1dc == EXMEMALUOut[9:0] ? DMemory_476 : _GEN_3704; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3706 = 10'h1dd == EXMEMALUOut[9:0] ? DMemory_477 : _GEN_3705; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3707 = 10'h1de == EXMEMALUOut[9:0] ? DMemory_478 : _GEN_3706; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3708 = 10'h1df == EXMEMALUOut[9:0] ? DMemory_479 : _GEN_3707; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3709 = 10'h1e0 == EXMEMALUOut[9:0] ? DMemory_480 : _GEN_3708; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3710 = 10'h1e1 == EXMEMALUOut[9:0] ? DMemory_481 : _GEN_3709; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3711 = 10'h1e2 == EXMEMALUOut[9:0] ? DMemory_482 : _GEN_3710; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3712 = 10'h1e3 == EXMEMALUOut[9:0] ? DMemory_483 : _GEN_3711; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3713 = 10'h1e4 == EXMEMALUOut[9:0] ? DMemory_484 : _GEN_3712; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3714 = 10'h1e5 == EXMEMALUOut[9:0] ? DMemory_485 : _GEN_3713; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3715 = 10'h1e6 == EXMEMALUOut[9:0] ? DMemory_486 : _GEN_3714; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3716 = 10'h1e7 == EXMEMALUOut[9:0] ? DMemory_487 : _GEN_3715; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3717 = 10'h1e8 == EXMEMALUOut[9:0] ? DMemory_488 : _GEN_3716; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3718 = 10'h1e9 == EXMEMALUOut[9:0] ? DMemory_489 : _GEN_3717; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3719 = 10'h1ea == EXMEMALUOut[9:0] ? DMemory_490 : _GEN_3718; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3720 = 10'h1eb == EXMEMALUOut[9:0] ? DMemory_491 : _GEN_3719; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3721 = 10'h1ec == EXMEMALUOut[9:0] ? DMemory_492 : _GEN_3720; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3722 = 10'h1ed == EXMEMALUOut[9:0] ? DMemory_493 : _GEN_3721; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3723 = 10'h1ee == EXMEMALUOut[9:0] ? DMemory_494 : _GEN_3722; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3724 = 10'h1ef == EXMEMALUOut[9:0] ? DMemory_495 : _GEN_3723; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3725 = 10'h1f0 == EXMEMALUOut[9:0] ? DMemory_496 : _GEN_3724; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3726 = 10'h1f1 == EXMEMALUOut[9:0] ? DMemory_497 : _GEN_3725; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3727 = 10'h1f2 == EXMEMALUOut[9:0] ? DMemory_498 : _GEN_3726; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3728 = 10'h1f3 == EXMEMALUOut[9:0] ? DMemory_499 : _GEN_3727; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3729 = 10'h1f4 == EXMEMALUOut[9:0] ? DMemory_500 : _GEN_3728; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3730 = 10'h1f5 == EXMEMALUOut[9:0] ? DMemory_501 : _GEN_3729; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3731 = 10'h1f6 == EXMEMALUOut[9:0] ? DMemory_502 : _GEN_3730; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3732 = 10'h1f7 == EXMEMALUOut[9:0] ? DMemory_503 : _GEN_3731; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3733 = 10'h1f8 == EXMEMALUOut[9:0] ? DMemory_504 : _GEN_3732; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3734 = 10'h1f9 == EXMEMALUOut[9:0] ? DMemory_505 : _GEN_3733; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3735 = 10'h1fa == EXMEMALUOut[9:0] ? DMemory_506 : _GEN_3734; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3736 = 10'h1fb == EXMEMALUOut[9:0] ? DMemory_507 : _GEN_3735; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3737 = 10'h1fc == EXMEMALUOut[9:0] ? DMemory_508 : _GEN_3736; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3738 = 10'h1fd == EXMEMALUOut[9:0] ? DMemory_509 : _GEN_3737; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3739 = 10'h1fe == EXMEMALUOut[9:0] ? DMemory_510 : _GEN_3738; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3740 = 10'h1ff == EXMEMALUOut[9:0] ? DMemory_511 : _GEN_3739; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3741 = 10'h200 == EXMEMALUOut[9:0] ? DMemory_512 : _GEN_3740; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3742 = 10'h201 == EXMEMALUOut[9:0] ? DMemory_513 : _GEN_3741; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3743 = 10'h202 == EXMEMALUOut[9:0] ? DMemory_514 : _GEN_3742; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3744 = 10'h203 == EXMEMALUOut[9:0] ? DMemory_515 : _GEN_3743; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3745 = 10'h204 == EXMEMALUOut[9:0] ? DMemory_516 : _GEN_3744; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3746 = 10'h205 == EXMEMALUOut[9:0] ? DMemory_517 : _GEN_3745; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3747 = 10'h206 == EXMEMALUOut[9:0] ? DMemory_518 : _GEN_3746; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3748 = 10'h207 == EXMEMALUOut[9:0] ? DMemory_519 : _GEN_3747; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3749 = 10'h208 == EXMEMALUOut[9:0] ? DMemory_520 : _GEN_3748; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3750 = 10'h209 == EXMEMALUOut[9:0] ? DMemory_521 : _GEN_3749; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3751 = 10'h20a == EXMEMALUOut[9:0] ? DMemory_522 : _GEN_3750; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3752 = 10'h20b == EXMEMALUOut[9:0] ? DMemory_523 : _GEN_3751; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3753 = 10'h20c == EXMEMALUOut[9:0] ? DMemory_524 : _GEN_3752; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3754 = 10'h20d == EXMEMALUOut[9:0] ? DMemory_525 : _GEN_3753; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3755 = 10'h20e == EXMEMALUOut[9:0] ? DMemory_526 : _GEN_3754; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3756 = 10'h20f == EXMEMALUOut[9:0] ? DMemory_527 : _GEN_3755; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3757 = 10'h210 == EXMEMALUOut[9:0] ? DMemory_528 : _GEN_3756; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3758 = 10'h211 == EXMEMALUOut[9:0] ? DMemory_529 : _GEN_3757; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3759 = 10'h212 == EXMEMALUOut[9:0] ? DMemory_530 : _GEN_3758; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3760 = 10'h213 == EXMEMALUOut[9:0] ? DMemory_531 : _GEN_3759; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3761 = 10'h214 == EXMEMALUOut[9:0] ? DMemory_532 : _GEN_3760; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3762 = 10'h215 == EXMEMALUOut[9:0] ? DMemory_533 : _GEN_3761; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3763 = 10'h216 == EXMEMALUOut[9:0] ? DMemory_534 : _GEN_3762; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3764 = 10'h217 == EXMEMALUOut[9:0] ? DMemory_535 : _GEN_3763; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3765 = 10'h218 == EXMEMALUOut[9:0] ? DMemory_536 : _GEN_3764; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3766 = 10'h219 == EXMEMALUOut[9:0] ? DMemory_537 : _GEN_3765; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3767 = 10'h21a == EXMEMALUOut[9:0] ? DMemory_538 : _GEN_3766; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3768 = 10'h21b == EXMEMALUOut[9:0] ? DMemory_539 : _GEN_3767; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3769 = 10'h21c == EXMEMALUOut[9:0] ? DMemory_540 : _GEN_3768; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3770 = 10'h21d == EXMEMALUOut[9:0] ? DMemory_541 : _GEN_3769; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3771 = 10'h21e == EXMEMALUOut[9:0] ? DMemory_542 : _GEN_3770; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3772 = 10'h21f == EXMEMALUOut[9:0] ? DMemory_543 : _GEN_3771; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3773 = 10'h220 == EXMEMALUOut[9:0] ? DMemory_544 : _GEN_3772; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3774 = 10'h221 == EXMEMALUOut[9:0] ? DMemory_545 : _GEN_3773; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3775 = 10'h222 == EXMEMALUOut[9:0] ? DMemory_546 : _GEN_3774; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3776 = 10'h223 == EXMEMALUOut[9:0] ? DMemory_547 : _GEN_3775; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3777 = 10'h224 == EXMEMALUOut[9:0] ? DMemory_548 : _GEN_3776; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3778 = 10'h225 == EXMEMALUOut[9:0] ? DMemory_549 : _GEN_3777; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3779 = 10'h226 == EXMEMALUOut[9:0] ? DMemory_550 : _GEN_3778; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3780 = 10'h227 == EXMEMALUOut[9:0] ? DMemory_551 : _GEN_3779; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3781 = 10'h228 == EXMEMALUOut[9:0] ? DMemory_552 : _GEN_3780; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3782 = 10'h229 == EXMEMALUOut[9:0] ? DMemory_553 : _GEN_3781; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3783 = 10'h22a == EXMEMALUOut[9:0] ? DMemory_554 : _GEN_3782; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3784 = 10'h22b == EXMEMALUOut[9:0] ? DMemory_555 : _GEN_3783; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3785 = 10'h22c == EXMEMALUOut[9:0] ? DMemory_556 : _GEN_3784; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3786 = 10'h22d == EXMEMALUOut[9:0] ? DMemory_557 : _GEN_3785; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3787 = 10'h22e == EXMEMALUOut[9:0] ? DMemory_558 : _GEN_3786; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3788 = 10'h22f == EXMEMALUOut[9:0] ? DMemory_559 : _GEN_3787; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3789 = 10'h230 == EXMEMALUOut[9:0] ? DMemory_560 : _GEN_3788; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3790 = 10'h231 == EXMEMALUOut[9:0] ? DMemory_561 : _GEN_3789; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3791 = 10'h232 == EXMEMALUOut[9:0] ? DMemory_562 : _GEN_3790; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3792 = 10'h233 == EXMEMALUOut[9:0] ? DMemory_563 : _GEN_3791; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3793 = 10'h234 == EXMEMALUOut[9:0] ? DMemory_564 : _GEN_3792; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3794 = 10'h235 == EXMEMALUOut[9:0] ? DMemory_565 : _GEN_3793; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3795 = 10'h236 == EXMEMALUOut[9:0] ? DMemory_566 : _GEN_3794; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3796 = 10'h237 == EXMEMALUOut[9:0] ? DMemory_567 : _GEN_3795; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3797 = 10'h238 == EXMEMALUOut[9:0] ? DMemory_568 : _GEN_3796; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3798 = 10'h239 == EXMEMALUOut[9:0] ? DMemory_569 : _GEN_3797; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3799 = 10'h23a == EXMEMALUOut[9:0] ? DMemory_570 : _GEN_3798; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3800 = 10'h23b == EXMEMALUOut[9:0] ? DMemory_571 : _GEN_3799; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3801 = 10'h23c == EXMEMALUOut[9:0] ? DMemory_572 : _GEN_3800; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3802 = 10'h23d == EXMEMALUOut[9:0] ? DMemory_573 : _GEN_3801; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3803 = 10'h23e == EXMEMALUOut[9:0] ? DMemory_574 : _GEN_3802; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3804 = 10'h23f == EXMEMALUOut[9:0] ? DMemory_575 : _GEN_3803; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3805 = 10'h240 == EXMEMALUOut[9:0] ? DMemory_576 : _GEN_3804; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3806 = 10'h241 == EXMEMALUOut[9:0] ? DMemory_577 : _GEN_3805; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3807 = 10'h242 == EXMEMALUOut[9:0] ? DMemory_578 : _GEN_3806; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3808 = 10'h243 == EXMEMALUOut[9:0] ? DMemory_579 : _GEN_3807; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3809 = 10'h244 == EXMEMALUOut[9:0] ? DMemory_580 : _GEN_3808; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3810 = 10'h245 == EXMEMALUOut[9:0] ? DMemory_581 : _GEN_3809; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3811 = 10'h246 == EXMEMALUOut[9:0] ? DMemory_582 : _GEN_3810; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3812 = 10'h247 == EXMEMALUOut[9:0] ? DMemory_583 : _GEN_3811; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3813 = 10'h248 == EXMEMALUOut[9:0] ? DMemory_584 : _GEN_3812; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3814 = 10'h249 == EXMEMALUOut[9:0] ? DMemory_585 : _GEN_3813; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3815 = 10'h24a == EXMEMALUOut[9:0] ? DMemory_586 : _GEN_3814; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3816 = 10'h24b == EXMEMALUOut[9:0] ? DMemory_587 : _GEN_3815; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3817 = 10'h24c == EXMEMALUOut[9:0] ? DMemory_588 : _GEN_3816; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3818 = 10'h24d == EXMEMALUOut[9:0] ? DMemory_589 : _GEN_3817; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3819 = 10'h24e == EXMEMALUOut[9:0] ? DMemory_590 : _GEN_3818; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3820 = 10'h24f == EXMEMALUOut[9:0] ? DMemory_591 : _GEN_3819; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3821 = 10'h250 == EXMEMALUOut[9:0] ? DMemory_592 : _GEN_3820; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3822 = 10'h251 == EXMEMALUOut[9:0] ? DMemory_593 : _GEN_3821; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3823 = 10'h252 == EXMEMALUOut[9:0] ? DMemory_594 : _GEN_3822; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3824 = 10'h253 == EXMEMALUOut[9:0] ? DMemory_595 : _GEN_3823; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3825 = 10'h254 == EXMEMALUOut[9:0] ? DMemory_596 : _GEN_3824; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3826 = 10'h255 == EXMEMALUOut[9:0] ? DMemory_597 : _GEN_3825; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3827 = 10'h256 == EXMEMALUOut[9:0] ? DMemory_598 : _GEN_3826; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3828 = 10'h257 == EXMEMALUOut[9:0] ? DMemory_599 : _GEN_3827; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3829 = 10'h258 == EXMEMALUOut[9:0] ? DMemory_600 : _GEN_3828; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3830 = 10'h259 == EXMEMALUOut[9:0] ? DMemory_601 : _GEN_3829; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3831 = 10'h25a == EXMEMALUOut[9:0] ? DMemory_602 : _GEN_3830; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3832 = 10'h25b == EXMEMALUOut[9:0] ? DMemory_603 : _GEN_3831; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3833 = 10'h25c == EXMEMALUOut[9:0] ? DMemory_604 : _GEN_3832; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3834 = 10'h25d == EXMEMALUOut[9:0] ? DMemory_605 : _GEN_3833; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3835 = 10'h25e == EXMEMALUOut[9:0] ? DMemory_606 : _GEN_3834; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3836 = 10'h25f == EXMEMALUOut[9:0] ? DMemory_607 : _GEN_3835; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3837 = 10'h260 == EXMEMALUOut[9:0] ? DMemory_608 : _GEN_3836; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3838 = 10'h261 == EXMEMALUOut[9:0] ? DMemory_609 : _GEN_3837; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3839 = 10'h262 == EXMEMALUOut[9:0] ? DMemory_610 : _GEN_3838; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3840 = 10'h263 == EXMEMALUOut[9:0] ? DMemory_611 : _GEN_3839; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3841 = 10'h264 == EXMEMALUOut[9:0] ? DMemory_612 : _GEN_3840; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3842 = 10'h265 == EXMEMALUOut[9:0] ? DMemory_613 : _GEN_3841; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3843 = 10'h266 == EXMEMALUOut[9:0] ? DMemory_614 : _GEN_3842; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3844 = 10'h267 == EXMEMALUOut[9:0] ? DMemory_615 : _GEN_3843; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3845 = 10'h268 == EXMEMALUOut[9:0] ? DMemory_616 : _GEN_3844; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3846 = 10'h269 == EXMEMALUOut[9:0] ? DMemory_617 : _GEN_3845; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3847 = 10'h26a == EXMEMALUOut[9:0] ? DMemory_618 : _GEN_3846; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3848 = 10'h26b == EXMEMALUOut[9:0] ? DMemory_619 : _GEN_3847; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3849 = 10'h26c == EXMEMALUOut[9:0] ? DMemory_620 : _GEN_3848; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3850 = 10'h26d == EXMEMALUOut[9:0] ? DMemory_621 : _GEN_3849; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3851 = 10'h26e == EXMEMALUOut[9:0] ? DMemory_622 : _GEN_3850; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3852 = 10'h26f == EXMEMALUOut[9:0] ? DMemory_623 : _GEN_3851; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3853 = 10'h270 == EXMEMALUOut[9:0] ? DMemory_624 : _GEN_3852; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3854 = 10'h271 == EXMEMALUOut[9:0] ? DMemory_625 : _GEN_3853; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3855 = 10'h272 == EXMEMALUOut[9:0] ? DMemory_626 : _GEN_3854; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3856 = 10'h273 == EXMEMALUOut[9:0] ? DMemory_627 : _GEN_3855; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3857 = 10'h274 == EXMEMALUOut[9:0] ? DMemory_628 : _GEN_3856; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3858 = 10'h275 == EXMEMALUOut[9:0] ? DMemory_629 : _GEN_3857; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3859 = 10'h276 == EXMEMALUOut[9:0] ? DMemory_630 : _GEN_3858; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3860 = 10'h277 == EXMEMALUOut[9:0] ? DMemory_631 : _GEN_3859; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3861 = 10'h278 == EXMEMALUOut[9:0] ? DMemory_632 : _GEN_3860; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3862 = 10'h279 == EXMEMALUOut[9:0] ? DMemory_633 : _GEN_3861; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3863 = 10'h27a == EXMEMALUOut[9:0] ? DMemory_634 : _GEN_3862; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3864 = 10'h27b == EXMEMALUOut[9:0] ? DMemory_635 : _GEN_3863; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3865 = 10'h27c == EXMEMALUOut[9:0] ? DMemory_636 : _GEN_3864; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3866 = 10'h27d == EXMEMALUOut[9:0] ? DMemory_637 : _GEN_3865; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3867 = 10'h27e == EXMEMALUOut[9:0] ? DMemory_638 : _GEN_3866; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3868 = 10'h27f == EXMEMALUOut[9:0] ? DMemory_639 : _GEN_3867; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3869 = 10'h280 == EXMEMALUOut[9:0] ? DMemory_640 : _GEN_3868; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3870 = 10'h281 == EXMEMALUOut[9:0] ? DMemory_641 : _GEN_3869; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3871 = 10'h282 == EXMEMALUOut[9:0] ? DMemory_642 : _GEN_3870; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3872 = 10'h283 == EXMEMALUOut[9:0] ? DMemory_643 : _GEN_3871; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3873 = 10'h284 == EXMEMALUOut[9:0] ? DMemory_644 : _GEN_3872; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3874 = 10'h285 == EXMEMALUOut[9:0] ? DMemory_645 : _GEN_3873; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3875 = 10'h286 == EXMEMALUOut[9:0] ? DMemory_646 : _GEN_3874; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3876 = 10'h287 == EXMEMALUOut[9:0] ? DMemory_647 : _GEN_3875; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3877 = 10'h288 == EXMEMALUOut[9:0] ? DMemory_648 : _GEN_3876; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3878 = 10'h289 == EXMEMALUOut[9:0] ? DMemory_649 : _GEN_3877; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3879 = 10'h28a == EXMEMALUOut[9:0] ? DMemory_650 : _GEN_3878; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3880 = 10'h28b == EXMEMALUOut[9:0] ? DMemory_651 : _GEN_3879; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3881 = 10'h28c == EXMEMALUOut[9:0] ? DMemory_652 : _GEN_3880; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3882 = 10'h28d == EXMEMALUOut[9:0] ? DMemory_653 : _GEN_3881; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3883 = 10'h28e == EXMEMALUOut[9:0] ? DMemory_654 : _GEN_3882; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3884 = 10'h28f == EXMEMALUOut[9:0] ? DMemory_655 : _GEN_3883; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3885 = 10'h290 == EXMEMALUOut[9:0] ? DMemory_656 : _GEN_3884; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3886 = 10'h291 == EXMEMALUOut[9:0] ? DMemory_657 : _GEN_3885; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3887 = 10'h292 == EXMEMALUOut[9:0] ? DMemory_658 : _GEN_3886; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3888 = 10'h293 == EXMEMALUOut[9:0] ? DMemory_659 : _GEN_3887; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3889 = 10'h294 == EXMEMALUOut[9:0] ? DMemory_660 : _GEN_3888; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3890 = 10'h295 == EXMEMALUOut[9:0] ? DMemory_661 : _GEN_3889; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3891 = 10'h296 == EXMEMALUOut[9:0] ? DMemory_662 : _GEN_3890; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3892 = 10'h297 == EXMEMALUOut[9:0] ? DMemory_663 : _GEN_3891; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3893 = 10'h298 == EXMEMALUOut[9:0] ? DMemory_664 : _GEN_3892; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3894 = 10'h299 == EXMEMALUOut[9:0] ? DMemory_665 : _GEN_3893; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3895 = 10'h29a == EXMEMALUOut[9:0] ? DMemory_666 : _GEN_3894; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3896 = 10'h29b == EXMEMALUOut[9:0] ? DMemory_667 : _GEN_3895; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3897 = 10'h29c == EXMEMALUOut[9:0] ? DMemory_668 : _GEN_3896; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3898 = 10'h29d == EXMEMALUOut[9:0] ? DMemory_669 : _GEN_3897; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3899 = 10'h29e == EXMEMALUOut[9:0] ? DMemory_670 : _GEN_3898; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3900 = 10'h29f == EXMEMALUOut[9:0] ? DMemory_671 : _GEN_3899; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3901 = 10'h2a0 == EXMEMALUOut[9:0] ? DMemory_672 : _GEN_3900; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3902 = 10'h2a1 == EXMEMALUOut[9:0] ? DMemory_673 : _GEN_3901; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3903 = 10'h2a2 == EXMEMALUOut[9:0] ? DMemory_674 : _GEN_3902; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3904 = 10'h2a3 == EXMEMALUOut[9:0] ? DMemory_675 : _GEN_3903; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3905 = 10'h2a4 == EXMEMALUOut[9:0] ? DMemory_676 : _GEN_3904; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3906 = 10'h2a5 == EXMEMALUOut[9:0] ? DMemory_677 : _GEN_3905; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3907 = 10'h2a6 == EXMEMALUOut[9:0] ? DMemory_678 : _GEN_3906; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3908 = 10'h2a7 == EXMEMALUOut[9:0] ? DMemory_679 : _GEN_3907; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3909 = 10'h2a8 == EXMEMALUOut[9:0] ? DMemory_680 : _GEN_3908; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3910 = 10'h2a9 == EXMEMALUOut[9:0] ? DMemory_681 : _GEN_3909; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3911 = 10'h2aa == EXMEMALUOut[9:0] ? DMemory_682 : _GEN_3910; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3912 = 10'h2ab == EXMEMALUOut[9:0] ? DMemory_683 : _GEN_3911; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3913 = 10'h2ac == EXMEMALUOut[9:0] ? DMemory_684 : _GEN_3912; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3914 = 10'h2ad == EXMEMALUOut[9:0] ? DMemory_685 : _GEN_3913; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3915 = 10'h2ae == EXMEMALUOut[9:0] ? DMemory_686 : _GEN_3914; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3916 = 10'h2af == EXMEMALUOut[9:0] ? DMemory_687 : _GEN_3915; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3917 = 10'h2b0 == EXMEMALUOut[9:0] ? DMemory_688 : _GEN_3916; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3918 = 10'h2b1 == EXMEMALUOut[9:0] ? DMemory_689 : _GEN_3917; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3919 = 10'h2b2 == EXMEMALUOut[9:0] ? DMemory_690 : _GEN_3918; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3920 = 10'h2b3 == EXMEMALUOut[9:0] ? DMemory_691 : _GEN_3919; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3921 = 10'h2b4 == EXMEMALUOut[9:0] ? DMemory_692 : _GEN_3920; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3922 = 10'h2b5 == EXMEMALUOut[9:0] ? DMemory_693 : _GEN_3921; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3923 = 10'h2b6 == EXMEMALUOut[9:0] ? DMemory_694 : _GEN_3922; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3924 = 10'h2b7 == EXMEMALUOut[9:0] ? DMemory_695 : _GEN_3923; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3925 = 10'h2b8 == EXMEMALUOut[9:0] ? DMemory_696 : _GEN_3924; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3926 = 10'h2b9 == EXMEMALUOut[9:0] ? DMemory_697 : _GEN_3925; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3927 = 10'h2ba == EXMEMALUOut[9:0] ? DMemory_698 : _GEN_3926; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3928 = 10'h2bb == EXMEMALUOut[9:0] ? DMemory_699 : _GEN_3927; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3929 = 10'h2bc == EXMEMALUOut[9:0] ? DMemory_700 : _GEN_3928; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3930 = 10'h2bd == EXMEMALUOut[9:0] ? DMemory_701 : _GEN_3929; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3931 = 10'h2be == EXMEMALUOut[9:0] ? DMemory_702 : _GEN_3930; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3932 = 10'h2bf == EXMEMALUOut[9:0] ? DMemory_703 : _GEN_3931; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3933 = 10'h2c0 == EXMEMALUOut[9:0] ? DMemory_704 : _GEN_3932; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3934 = 10'h2c1 == EXMEMALUOut[9:0] ? DMemory_705 : _GEN_3933; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3935 = 10'h2c2 == EXMEMALUOut[9:0] ? DMemory_706 : _GEN_3934; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3936 = 10'h2c3 == EXMEMALUOut[9:0] ? DMemory_707 : _GEN_3935; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3937 = 10'h2c4 == EXMEMALUOut[9:0] ? DMemory_708 : _GEN_3936; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3938 = 10'h2c5 == EXMEMALUOut[9:0] ? DMemory_709 : _GEN_3937; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3939 = 10'h2c6 == EXMEMALUOut[9:0] ? DMemory_710 : _GEN_3938; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3940 = 10'h2c7 == EXMEMALUOut[9:0] ? DMemory_711 : _GEN_3939; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3941 = 10'h2c8 == EXMEMALUOut[9:0] ? DMemory_712 : _GEN_3940; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3942 = 10'h2c9 == EXMEMALUOut[9:0] ? DMemory_713 : _GEN_3941; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3943 = 10'h2ca == EXMEMALUOut[9:0] ? DMemory_714 : _GEN_3942; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3944 = 10'h2cb == EXMEMALUOut[9:0] ? DMemory_715 : _GEN_3943; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3945 = 10'h2cc == EXMEMALUOut[9:0] ? DMemory_716 : _GEN_3944; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3946 = 10'h2cd == EXMEMALUOut[9:0] ? DMemory_717 : _GEN_3945; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3947 = 10'h2ce == EXMEMALUOut[9:0] ? DMemory_718 : _GEN_3946; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3948 = 10'h2cf == EXMEMALUOut[9:0] ? DMemory_719 : _GEN_3947; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3949 = 10'h2d0 == EXMEMALUOut[9:0] ? DMemory_720 : _GEN_3948; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3950 = 10'h2d1 == EXMEMALUOut[9:0] ? DMemory_721 : _GEN_3949; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3951 = 10'h2d2 == EXMEMALUOut[9:0] ? DMemory_722 : _GEN_3950; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3952 = 10'h2d3 == EXMEMALUOut[9:0] ? DMemory_723 : _GEN_3951; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3953 = 10'h2d4 == EXMEMALUOut[9:0] ? DMemory_724 : _GEN_3952; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3954 = 10'h2d5 == EXMEMALUOut[9:0] ? DMemory_725 : _GEN_3953; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3955 = 10'h2d6 == EXMEMALUOut[9:0] ? DMemory_726 : _GEN_3954; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3956 = 10'h2d7 == EXMEMALUOut[9:0] ? DMemory_727 : _GEN_3955; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3957 = 10'h2d8 == EXMEMALUOut[9:0] ? DMemory_728 : _GEN_3956; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3958 = 10'h2d9 == EXMEMALUOut[9:0] ? DMemory_729 : _GEN_3957; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3959 = 10'h2da == EXMEMALUOut[9:0] ? DMemory_730 : _GEN_3958; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3960 = 10'h2db == EXMEMALUOut[9:0] ? DMemory_731 : _GEN_3959; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3961 = 10'h2dc == EXMEMALUOut[9:0] ? DMemory_732 : _GEN_3960; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3962 = 10'h2dd == EXMEMALUOut[9:0] ? DMemory_733 : _GEN_3961; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3963 = 10'h2de == EXMEMALUOut[9:0] ? DMemory_734 : _GEN_3962; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3964 = 10'h2df == EXMEMALUOut[9:0] ? DMemory_735 : _GEN_3963; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3965 = 10'h2e0 == EXMEMALUOut[9:0] ? DMemory_736 : _GEN_3964; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3966 = 10'h2e1 == EXMEMALUOut[9:0] ? DMemory_737 : _GEN_3965; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3967 = 10'h2e2 == EXMEMALUOut[9:0] ? DMemory_738 : _GEN_3966; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3968 = 10'h2e3 == EXMEMALUOut[9:0] ? DMemory_739 : _GEN_3967; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3969 = 10'h2e4 == EXMEMALUOut[9:0] ? DMemory_740 : _GEN_3968; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3970 = 10'h2e5 == EXMEMALUOut[9:0] ? DMemory_741 : _GEN_3969; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3971 = 10'h2e6 == EXMEMALUOut[9:0] ? DMemory_742 : _GEN_3970; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3972 = 10'h2e7 == EXMEMALUOut[9:0] ? DMemory_743 : _GEN_3971; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3973 = 10'h2e8 == EXMEMALUOut[9:0] ? DMemory_744 : _GEN_3972; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3974 = 10'h2e9 == EXMEMALUOut[9:0] ? DMemory_745 : _GEN_3973; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3975 = 10'h2ea == EXMEMALUOut[9:0] ? DMemory_746 : _GEN_3974; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3976 = 10'h2eb == EXMEMALUOut[9:0] ? DMemory_747 : _GEN_3975; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3977 = 10'h2ec == EXMEMALUOut[9:0] ? DMemory_748 : _GEN_3976; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3978 = 10'h2ed == EXMEMALUOut[9:0] ? DMemory_749 : _GEN_3977; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3979 = 10'h2ee == EXMEMALUOut[9:0] ? DMemory_750 : _GEN_3978; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3980 = 10'h2ef == EXMEMALUOut[9:0] ? DMemory_751 : _GEN_3979; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3981 = 10'h2f0 == EXMEMALUOut[9:0] ? DMemory_752 : _GEN_3980; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3982 = 10'h2f1 == EXMEMALUOut[9:0] ? DMemory_753 : _GEN_3981; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3983 = 10'h2f2 == EXMEMALUOut[9:0] ? DMemory_754 : _GEN_3982; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3984 = 10'h2f3 == EXMEMALUOut[9:0] ? DMemory_755 : _GEN_3983; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3985 = 10'h2f4 == EXMEMALUOut[9:0] ? DMemory_756 : _GEN_3984; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3986 = 10'h2f5 == EXMEMALUOut[9:0] ? DMemory_757 : _GEN_3985; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3987 = 10'h2f6 == EXMEMALUOut[9:0] ? DMemory_758 : _GEN_3986; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3988 = 10'h2f7 == EXMEMALUOut[9:0] ? DMemory_759 : _GEN_3987; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3989 = 10'h2f8 == EXMEMALUOut[9:0] ? DMemory_760 : _GEN_3988; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3990 = 10'h2f9 == EXMEMALUOut[9:0] ? DMemory_761 : _GEN_3989; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3991 = 10'h2fa == EXMEMALUOut[9:0] ? DMemory_762 : _GEN_3990; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3992 = 10'h2fb == EXMEMALUOut[9:0] ? DMemory_763 : _GEN_3991; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3993 = 10'h2fc == EXMEMALUOut[9:0] ? DMemory_764 : _GEN_3992; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3994 = 10'h2fd == EXMEMALUOut[9:0] ? DMemory_765 : _GEN_3993; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3995 = 10'h2fe == EXMEMALUOut[9:0] ? DMemory_766 : _GEN_3994; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3996 = 10'h2ff == EXMEMALUOut[9:0] ? DMemory_767 : _GEN_3995; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3997 = 10'h300 == EXMEMALUOut[9:0] ? DMemory_768 : _GEN_3996; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3998 = 10'h301 == EXMEMALUOut[9:0] ? DMemory_769 : _GEN_3997; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_3999 = 10'h302 == EXMEMALUOut[9:0] ? DMemory_770 : _GEN_3998; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4000 = 10'h303 == EXMEMALUOut[9:0] ? DMemory_771 : _GEN_3999; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4001 = 10'h304 == EXMEMALUOut[9:0] ? DMemory_772 : _GEN_4000; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4002 = 10'h305 == EXMEMALUOut[9:0] ? DMemory_773 : _GEN_4001; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4003 = 10'h306 == EXMEMALUOut[9:0] ? DMemory_774 : _GEN_4002; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4004 = 10'h307 == EXMEMALUOut[9:0] ? DMemory_775 : _GEN_4003; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4005 = 10'h308 == EXMEMALUOut[9:0] ? DMemory_776 : _GEN_4004; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4006 = 10'h309 == EXMEMALUOut[9:0] ? DMemory_777 : _GEN_4005; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4007 = 10'h30a == EXMEMALUOut[9:0] ? DMemory_778 : _GEN_4006; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4008 = 10'h30b == EXMEMALUOut[9:0] ? DMemory_779 : _GEN_4007; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4009 = 10'h30c == EXMEMALUOut[9:0] ? DMemory_780 : _GEN_4008; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4010 = 10'h30d == EXMEMALUOut[9:0] ? DMemory_781 : _GEN_4009; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4011 = 10'h30e == EXMEMALUOut[9:0] ? DMemory_782 : _GEN_4010; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4012 = 10'h30f == EXMEMALUOut[9:0] ? DMemory_783 : _GEN_4011; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4013 = 10'h310 == EXMEMALUOut[9:0] ? DMemory_784 : _GEN_4012; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4014 = 10'h311 == EXMEMALUOut[9:0] ? DMemory_785 : _GEN_4013; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4015 = 10'h312 == EXMEMALUOut[9:0] ? DMemory_786 : _GEN_4014; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4016 = 10'h313 == EXMEMALUOut[9:0] ? DMemory_787 : _GEN_4015; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4017 = 10'h314 == EXMEMALUOut[9:0] ? DMemory_788 : _GEN_4016; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4018 = 10'h315 == EXMEMALUOut[9:0] ? DMemory_789 : _GEN_4017; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4019 = 10'h316 == EXMEMALUOut[9:0] ? DMemory_790 : _GEN_4018; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4020 = 10'h317 == EXMEMALUOut[9:0] ? DMemory_791 : _GEN_4019; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4021 = 10'h318 == EXMEMALUOut[9:0] ? DMemory_792 : _GEN_4020; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4022 = 10'h319 == EXMEMALUOut[9:0] ? DMemory_793 : _GEN_4021; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4023 = 10'h31a == EXMEMALUOut[9:0] ? DMemory_794 : _GEN_4022; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4024 = 10'h31b == EXMEMALUOut[9:0] ? DMemory_795 : _GEN_4023; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4025 = 10'h31c == EXMEMALUOut[9:0] ? DMemory_796 : _GEN_4024; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4026 = 10'h31d == EXMEMALUOut[9:0] ? DMemory_797 : _GEN_4025; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4027 = 10'h31e == EXMEMALUOut[9:0] ? DMemory_798 : _GEN_4026; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4028 = 10'h31f == EXMEMALUOut[9:0] ? DMemory_799 : _GEN_4027; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4029 = 10'h320 == EXMEMALUOut[9:0] ? DMemory_800 : _GEN_4028; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4030 = 10'h321 == EXMEMALUOut[9:0] ? DMemory_801 : _GEN_4029; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4031 = 10'h322 == EXMEMALUOut[9:0] ? DMemory_802 : _GEN_4030; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4032 = 10'h323 == EXMEMALUOut[9:0] ? DMemory_803 : _GEN_4031; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4033 = 10'h324 == EXMEMALUOut[9:0] ? DMemory_804 : _GEN_4032; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4034 = 10'h325 == EXMEMALUOut[9:0] ? DMemory_805 : _GEN_4033; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4035 = 10'h326 == EXMEMALUOut[9:0] ? DMemory_806 : _GEN_4034; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4036 = 10'h327 == EXMEMALUOut[9:0] ? DMemory_807 : _GEN_4035; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4037 = 10'h328 == EXMEMALUOut[9:0] ? DMemory_808 : _GEN_4036; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4038 = 10'h329 == EXMEMALUOut[9:0] ? DMemory_809 : _GEN_4037; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4039 = 10'h32a == EXMEMALUOut[9:0] ? DMemory_810 : _GEN_4038; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4040 = 10'h32b == EXMEMALUOut[9:0] ? DMemory_811 : _GEN_4039; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4041 = 10'h32c == EXMEMALUOut[9:0] ? DMemory_812 : _GEN_4040; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4042 = 10'h32d == EXMEMALUOut[9:0] ? DMemory_813 : _GEN_4041; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4043 = 10'h32e == EXMEMALUOut[9:0] ? DMemory_814 : _GEN_4042; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4044 = 10'h32f == EXMEMALUOut[9:0] ? DMemory_815 : _GEN_4043; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4045 = 10'h330 == EXMEMALUOut[9:0] ? DMemory_816 : _GEN_4044; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4046 = 10'h331 == EXMEMALUOut[9:0] ? DMemory_817 : _GEN_4045; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4047 = 10'h332 == EXMEMALUOut[9:0] ? DMemory_818 : _GEN_4046; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4048 = 10'h333 == EXMEMALUOut[9:0] ? DMemory_819 : _GEN_4047; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4049 = 10'h334 == EXMEMALUOut[9:0] ? DMemory_820 : _GEN_4048; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4050 = 10'h335 == EXMEMALUOut[9:0] ? DMemory_821 : _GEN_4049; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4051 = 10'h336 == EXMEMALUOut[9:0] ? DMemory_822 : _GEN_4050; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4052 = 10'h337 == EXMEMALUOut[9:0] ? DMemory_823 : _GEN_4051; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4053 = 10'h338 == EXMEMALUOut[9:0] ? DMemory_824 : _GEN_4052; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4054 = 10'h339 == EXMEMALUOut[9:0] ? DMemory_825 : _GEN_4053; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4055 = 10'h33a == EXMEMALUOut[9:0] ? DMemory_826 : _GEN_4054; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4056 = 10'h33b == EXMEMALUOut[9:0] ? DMemory_827 : _GEN_4055; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4057 = 10'h33c == EXMEMALUOut[9:0] ? DMemory_828 : _GEN_4056; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4058 = 10'h33d == EXMEMALUOut[9:0] ? DMemory_829 : _GEN_4057; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4059 = 10'h33e == EXMEMALUOut[9:0] ? DMemory_830 : _GEN_4058; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4060 = 10'h33f == EXMEMALUOut[9:0] ? DMemory_831 : _GEN_4059; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4061 = 10'h340 == EXMEMALUOut[9:0] ? DMemory_832 : _GEN_4060; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4062 = 10'h341 == EXMEMALUOut[9:0] ? DMemory_833 : _GEN_4061; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4063 = 10'h342 == EXMEMALUOut[9:0] ? DMemory_834 : _GEN_4062; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4064 = 10'h343 == EXMEMALUOut[9:0] ? DMemory_835 : _GEN_4063; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4065 = 10'h344 == EXMEMALUOut[9:0] ? DMemory_836 : _GEN_4064; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4066 = 10'h345 == EXMEMALUOut[9:0] ? DMemory_837 : _GEN_4065; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4067 = 10'h346 == EXMEMALUOut[9:0] ? DMemory_838 : _GEN_4066; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4068 = 10'h347 == EXMEMALUOut[9:0] ? DMemory_839 : _GEN_4067; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4069 = 10'h348 == EXMEMALUOut[9:0] ? DMemory_840 : _GEN_4068; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4070 = 10'h349 == EXMEMALUOut[9:0] ? DMemory_841 : _GEN_4069; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4071 = 10'h34a == EXMEMALUOut[9:0] ? DMemory_842 : _GEN_4070; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4072 = 10'h34b == EXMEMALUOut[9:0] ? DMemory_843 : _GEN_4071; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4073 = 10'h34c == EXMEMALUOut[9:0] ? DMemory_844 : _GEN_4072; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4074 = 10'h34d == EXMEMALUOut[9:0] ? DMemory_845 : _GEN_4073; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4075 = 10'h34e == EXMEMALUOut[9:0] ? DMemory_846 : _GEN_4074; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4076 = 10'h34f == EXMEMALUOut[9:0] ? DMemory_847 : _GEN_4075; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4077 = 10'h350 == EXMEMALUOut[9:0] ? DMemory_848 : _GEN_4076; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4078 = 10'h351 == EXMEMALUOut[9:0] ? DMemory_849 : _GEN_4077; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4079 = 10'h352 == EXMEMALUOut[9:0] ? DMemory_850 : _GEN_4078; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4080 = 10'h353 == EXMEMALUOut[9:0] ? DMemory_851 : _GEN_4079; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4081 = 10'h354 == EXMEMALUOut[9:0] ? DMemory_852 : _GEN_4080; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4082 = 10'h355 == EXMEMALUOut[9:0] ? DMemory_853 : _GEN_4081; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4083 = 10'h356 == EXMEMALUOut[9:0] ? DMemory_854 : _GEN_4082; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4084 = 10'h357 == EXMEMALUOut[9:0] ? DMemory_855 : _GEN_4083; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4085 = 10'h358 == EXMEMALUOut[9:0] ? DMemory_856 : _GEN_4084; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4086 = 10'h359 == EXMEMALUOut[9:0] ? DMemory_857 : _GEN_4085; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4087 = 10'h35a == EXMEMALUOut[9:0] ? DMemory_858 : _GEN_4086; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4088 = 10'h35b == EXMEMALUOut[9:0] ? DMemory_859 : _GEN_4087; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4089 = 10'h35c == EXMEMALUOut[9:0] ? DMemory_860 : _GEN_4088; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4090 = 10'h35d == EXMEMALUOut[9:0] ? DMemory_861 : _GEN_4089; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4091 = 10'h35e == EXMEMALUOut[9:0] ? DMemory_862 : _GEN_4090; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4092 = 10'h35f == EXMEMALUOut[9:0] ? DMemory_863 : _GEN_4091; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4093 = 10'h360 == EXMEMALUOut[9:0] ? DMemory_864 : _GEN_4092; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4094 = 10'h361 == EXMEMALUOut[9:0] ? DMemory_865 : _GEN_4093; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4095 = 10'h362 == EXMEMALUOut[9:0] ? DMemory_866 : _GEN_4094; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4096 = 10'h363 == EXMEMALUOut[9:0] ? DMemory_867 : _GEN_4095; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4097 = 10'h364 == EXMEMALUOut[9:0] ? DMemory_868 : _GEN_4096; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4098 = 10'h365 == EXMEMALUOut[9:0] ? DMemory_869 : _GEN_4097; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4099 = 10'h366 == EXMEMALUOut[9:0] ? DMemory_870 : _GEN_4098; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4100 = 10'h367 == EXMEMALUOut[9:0] ? DMemory_871 : _GEN_4099; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4101 = 10'h368 == EXMEMALUOut[9:0] ? DMemory_872 : _GEN_4100; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4102 = 10'h369 == EXMEMALUOut[9:0] ? DMemory_873 : _GEN_4101; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4103 = 10'h36a == EXMEMALUOut[9:0] ? DMemory_874 : _GEN_4102; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4104 = 10'h36b == EXMEMALUOut[9:0] ? DMemory_875 : _GEN_4103; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4105 = 10'h36c == EXMEMALUOut[9:0] ? DMemory_876 : _GEN_4104; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4106 = 10'h36d == EXMEMALUOut[9:0] ? DMemory_877 : _GEN_4105; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4107 = 10'h36e == EXMEMALUOut[9:0] ? DMemory_878 : _GEN_4106; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4108 = 10'h36f == EXMEMALUOut[9:0] ? DMemory_879 : _GEN_4107; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4109 = 10'h370 == EXMEMALUOut[9:0] ? DMemory_880 : _GEN_4108; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4110 = 10'h371 == EXMEMALUOut[9:0] ? DMemory_881 : _GEN_4109; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4111 = 10'h372 == EXMEMALUOut[9:0] ? DMemory_882 : _GEN_4110; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4112 = 10'h373 == EXMEMALUOut[9:0] ? DMemory_883 : _GEN_4111; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4113 = 10'h374 == EXMEMALUOut[9:0] ? DMemory_884 : _GEN_4112; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4114 = 10'h375 == EXMEMALUOut[9:0] ? DMemory_885 : _GEN_4113; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4115 = 10'h376 == EXMEMALUOut[9:0] ? DMemory_886 : _GEN_4114; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4116 = 10'h377 == EXMEMALUOut[9:0] ? DMemory_887 : _GEN_4115; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4117 = 10'h378 == EXMEMALUOut[9:0] ? DMemory_888 : _GEN_4116; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4118 = 10'h379 == EXMEMALUOut[9:0] ? DMemory_889 : _GEN_4117; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4119 = 10'h37a == EXMEMALUOut[9:0] ? DMemory_890 : _GEN_4118; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4120 = 10'h37b == EXMEMALUOut[9:0] ? DMemory_891 : _GEN_4119; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4121 = 10'h37c == EXMEMALUOut[9:0] ? DMemory_892 : _GEN_4120; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4122 = 10'h37d == EXMEMALUOut[9:0] ? DMemory_893 : _GEN_4121; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4123 = 10'h37e == EXMEMALUOut[9:0] ? DMemory_894 : _GEN_4122; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4124 = 10'h37f == EXMEMALUOut[9:0] ? DMemory_895 : _GEN_4123; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4125 = 10'h380 == EXMEMALUOut[9:0] ? DMemory_896 : _GEN_4124; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4126 = 10'h381 == EXMEMALUOut[9:0] ? DMemory_897 : _GEN_4125; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4127 = 10'h382 == EXMEMALUOut[9:0] ? DMemory_898 : _GEN_4126; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4128 = 10'h383 == EXMEMALUOut[9:0] ? DMemory_899 : _GEN_4127; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4129 = 10'h384 == EXMEMALUOut[9:0] ? DMemory_900 : _GEN_4128; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4130 = 10'h385 == EXMEMALUOut[9:0] ? DMemory_901 : _GEN_4129; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4131 = 10'h386 == EXMEMALUOut[9:0] ? DMemory_902 : _GEN_4130; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4132 = 10'h387 == EXMEMALUOut[9:0] ? DMemory_903 : _GEN_4131; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4133 = 10'h388 == EXMEMALUOut[9:0] ? DMemory_904 : _GEN_4132; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4134 = 10'h389 == EXMEMALUOut[9:0] ? DMemory_905 : _GEN_4133; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4135 = 10'h38a == EXMEMALUOut[9:0] ? DMemory_906 : _GEN_4134; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4136 = 10'h38b == EXMEMALUOut[9:0] ? DMemory_907 : _GEN_4135; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4137 = 10'h38c == EXMEMALUOut[9:0] ? DMemory_908 : _GEN_4136; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4138 = 10'h38d == EXMEMALUOut[9:0] ? DMemory_909 : _GEN_4137; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4139 = 10'h38e == EXMEMALUOut[9:0] ? DMemory_910 : _GEN_4138; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4140 = 10'h38f == EXMEMALUOut[9:0] ? DMemory_911 : _GEN_4139; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4141 = 10'h390 == EXMEMALUOut[9:0] ? DMemory_912 : _GEN_4140; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4142 = 10'h391 == EXMEMALUOut[9:0] ? DMemory_913 : _GEN_4141; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4143 = 10'h392 == EXMEMALUOut[9:0] ? DMemory_914 : _GEN_4142; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4144 = 10'h393 == EXMEMALUOut[9:0] ? DMemory_915 : _GEN_4143; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4145 = 10'h394 == EXMEMALUOut[9:0] ? DMemory_916 : _GEN_4144; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4146 = 10'h395 == EXMEMALUOut[9:0] ? DMemory_917 : _GEN_4145; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4147 = 10'h396 == EXMEMALUOut[9:0] ? DMemory_918 : _GEN_4146; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4148 = 10'h397 == EXMEMALUOut[9:0] ? DMemory_919 : _GEN_4147; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4149 = 10'h398 == EXMEMALUOut[9:0] ? DMemory_920 : _GEN_4148; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4150 = 10'h399 == EXMEMALUOut[9:0] ? DMemory_921 : _GEN_4149; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4151 = 10'h39a == EXMEMALUOut[9:0] ? DMemory_922 : _GEN_4150; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4152 = 10'h39b == EXMEMALUOut[9:0] ? DMemory_923 : _GEN_4151; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4153 = 10'h39c == EXMEMALUOut[9:0] ? DMemory_924 : _GEN_4152; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4154 = 10'h39d == EXMEMALUOut[9:0] ? DMemory_925 : _GEN_4153; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4155 = 10'h39e == EXMEMALUOut[9:0] ? DMemory_926 : _GEN_4154; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4156 = 10'h39f == EXMEMALUOut[9:0] ? DMemory_927 : _GEN_4155; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4157 = 10'h3a0 == EXMEMALUOut[9:0] ? DMemory_928 : _GEN_4156; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4158 = 10'h3a1 == EXMEMALUOut[9:0] ? DMemory_929 : _GEN_4157; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4159 = 10'h3a2 == EXMEMALUOut[9:0] ? DMemory_930 : _GEN_4158; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4160 = 10'h3a3 == EXMEMALUOut[9:0] ? DMemory_931 : _GEN_4159; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4161 = 10'h3a4 == EXMEMALUOut[9:0] ? DMemory_932 : _GEN_4160; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4162 = 10'h3a5 == EXMEMALUOut[9:0] ? DMemory_933 : _GEN_4161; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4163 = 10'h3a6 == EXMEMALUOut[9:0] ? DMemory_934 : _GEN_4162; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4164 = 10'h3a7 == EXMEMALUOut[9:0] ? DMemory_935 : _GEN_4163; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4165 = 10'h3a8 == EXMEMALUOut[9:0] ? DMemory_936 : _GEN_4164; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4166 = 10'h3a9 == EXMEMALUOut[9:0] ? DMemory_937 : _GEN_4165; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4167 = 10'h3aa == EXMEMALUOut[9:0] ? DMemory_938 : _GEN_4166; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4168 = 10'h3ab == EXMEMALUOut[9:0] ? DMemory_939 : _GEN_4167; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4169 = 10'h3ac == EXMEMALUOut[9:0] ? DMemory_940 : _GEN_4168; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4170 = 10'h3ad == EXMEMALUOut[9:0] ? DMemory_941 : _GEN_4169; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4171 = 10'h3ae == EXMEMALUOut[9:0] ? DMemory_942 : _GEN_4170; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4172 = 10'h3af == EXMEMALUOut[9:0] ? DMemory_943 : _GEN_4171; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4173 = 10'h3b0 == EXMEMALUOut[9:0] ? DMemory_944 : _GEN_4172; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4174 = 10'h3b1 == EXMEMALUOut[9:0] ? DMemory_945 : _GEN_4173; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4175 = 10'h3b2 == EXMEMALUOut[9:0] ? DMemory_946 : _GEN_4174; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4176 = 10'h3b3 == EXMEMALUOut[9:0] ? DMemory_947 : _GEN_4175; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4177 = 10'h3b4 == EXMEMALUOut[9:0] ? DMemory_948 : _GEN_4176; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4178 = 10'h3b5 == EXMEMALUOut[9:0] ? DMemory_949 : _GEN_4177; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4179 = 10'h3b6 == EXMEMALUOut[9:0] ? DMemory_950 : _GEN_4178; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4180 = 10'h3b7 == EXMEMALUOut[9:0] ? DMemory_951 : _GEN_4179; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4181 = 10'h3b8 == EXMEMALUOut[9:0] ? DMemory_952 : _GEN_4180; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4182 = 10'h3b9 == EXMEMALUOut[9:0] ? DMemory_953 : _GEN_4181; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4183 = 10'h3ba == EXMEMALUOut[9:0] ? DMemory_954 : _GEN_4182; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4184 = 10'h3bb == EXMEMALUOut[9:0] ? DMemory_955 : _GEN_4183; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4185 = 10'h3bc == EXMEMALUOut[9:0] ? DMemory_956 : _GEN_4184; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4186 = 10'h3bd == EXMEMALUOut[9:0] ? DMemory_957 : _GEN_4185; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4187 = 10'h3be == EXMEMALUOut[9:0] ? DMemory_958 : _GEN_4186; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4188 = 10'h3bf == EXMEMALUOut[9:0] ? DMemory_959 : _GEN_4187; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4189 = 10'h3c0 == EXMEMALUOut[9:0] ? DMemory_960 : _GEN_4188; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4190 = 10'h3c1 == EXMEMALUOut[9:0] ? DMemory_961 : _GEN_4189; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4191 = 10'h3c2 == EXMEMALUOut[9:0] ? DMemory_962 : _GEN_4190; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4192 = 10'h3c3 == EXMEMALUOut[9:0] ? DMemory_963 : _GEN_4191; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4193 = 10'h3c4 == EXMEMALUOut[9:0] ? DMemory_964 : _GEN_4192; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4194 = 10'h3c5 == EXMEMALUOut[9:0] ? DMemory_965 : _GEN_4193; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4195 = 10'h3c6 == EXMEMALUOut[9:0] ? DMemory_966 : _GEN_4194; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4196 = 10'h3c7 == EXMEMALUOut[9:0] ? DMemory_967 : _GEN_4195; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4197 = 10'h3c8 == EXMEMALUOut[9:0] ? DMemory_968 : _GEN_4196; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4198 = 10'h3c9 == EXMEMALUOut[9:0] ? DMemory_969 : _GEN_4197; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4199 = 10'h3ca == EXMEMALUOut[9:0] ? DMemory_970 : _GEN_4198; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4200 = 10'h3cb == EXMEMALUOut[9:0] ? DMemory_971 : _GEN_4199; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4201 = 10'h3cc == EXMEMALUOut[9:0] ? DMemory_972 : _GEN_4200; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4202 = 10'h3cd == EXMEMALUOut[9:0] ? DMemory_973 : _GEN_4201; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4203 = 10'h3ce == EXMEMALUOut[9:0] ? DMemory_974 : _GEN_4202; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4204 = 10'h3cf == EXMEMALUOut[9:0] ? DMemory_975 : _GEN_4203; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4205 = 10'h3d0 == EXMEMALUOut[9:0] ? DMemory_976 : _GEN_4204; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4206 = 10'h3d1 == EXMEMALUOut[9:0] ? DMemory_977 : _GEN_4205; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4207 = 10'h3d2 == EXMEMALUOut[9:0] ? DMemory_978 : _GEN_4206; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4208 = 10'h3d3 == EXMEMALUOut[9:0] ? DMemory_979 : _GEN_4207; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4209 = 10'h3d4 == EXMEMALUOut[9:0] ? DMemory_980 : _GEN_4208; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4210 = 10'h3d5 == EXMEMALUOut[9:0] ? DMemory_981 : _GEN_4209; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4211 = 10'h3d6 == EXMEMALUOut[9:0] ? DMemory_982 : _GEN_4210; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4212 = 10'h3d7 == EXMEMALUOut[9:0] ? DMemory_983 : _GEN_4211; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4213 = 10'h3d8 == EXMEMALUOut[9:0] ? DMemory_984 : _GEN_4212; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4214 = 10'h3d9 == EXMEMALUOut[9:0] ? DMemory_985 : _GEN_4213; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4215 = 10'h3da == EXMEMALUOut[9:0] ? DMemory_986 : _GEN_4214; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4216 = 10'h3db == EXMEMALUOut[9:0] ? DMemory_987 : _GEN_4215; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4217 = 10'h3dc == EXMEMALUOut[9:0] ? DMemory_988 : _GEN_4216; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4218 = 10'h3dd == EXMEMALUOut[9:0] ? DMemory_989 : _GEN_4217; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4219 = 10'h3de == EXMEMALUOut[9:0] ? DMemory_990 : _GEN_4218; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4220 = 10'h3df == EXMEMALUOut[9:0] ? DMemory_991 : _GEN_4219; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4221 = 10'h3e0 == EXMEMALUOut[9:0] ? DMemory_992 : _GEN_4220; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4222 = 10'h3e1 == EXMEMALUOut[9:0] ? DMemory_993 : _GEN_4221; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4223 = 10'h3e2 == EXMEMALUOut[9:0] ? DMemory_994 : _GEN_4222; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4224 = 10'h3e3 == EXMEMALUOut[9:0] ? DMemory_995 : _GEN_4223; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4225 = 10'h3e4 == EXMEMALUOut[9:0] ? DMemory_996 : _GEN_4224; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4226 = 10'h3e5 == EXMEMALUOut[9:0] ? DMemory_997 : _GEN_4225; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4227 = 10'h3e6 == EXMEMALUOut[9:0] ? DMemory_998 : _GEN_4226; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4228 = 10'h3e7 == EXMEMALUOut[9:0] ? DMemory_999 : _GEN_4227; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4229 = 10'h3e8 == EXMEMALUOut[9:0] ? DMemory_1000 : _GEN_4228; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4230 = 10'h3e9 == EXMEMALUOut[9:0] ? DMemory_1001 : _GEN_4229; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4231 = 10'h3ea == EXMEMALUOut[9:0] ? DMemory_1002 : _GEN_4230; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4232 = 10'h3eb == EXMEMALUOut[9:0] ? DMemory_1003 : _GEN_4231; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4233 = 10'h3ec == EXMEMALUOut[9:0] ? DMemory_1004 : _GEN_4232; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4234 = 10'h3ed == EXMEMALUOut[9:0] ? DMemory_1005 : _GEN_4233; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4235 = 10'h3ee == EXMEMALUOut[9:0] ? DMemory_1006 : _GEN_4234; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4236 = 10'h3ef == EXMEMALUOut[9:0] ? DMemory_1007 : _GEN_4235; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4237 = 10'h3f0 == EXMEMALUOut[9:0] ? DMemory_1008 : _GEN_4236; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4238 = 10'h3f1 == EXMEMALUOut[9:0] ? DMemory_1009 : _GEN_4237; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4239 = 10'h3f2 == EXMEMALUOut[9:0] ? DMemory_1010 : _GEN_4238; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4240 = 10'h3f3 == EXMEMALUOut[9:0] ? DMemory_1011 : _GEN_4239; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4241 = 10'h3f4 == EXMEMALUOut[9:0] ? DMemory_1012 : _GEN_4240; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4242 = 10'h3f5 == EXMEMALUOut[9:0] ? DMemory_1013 : _GEN_4241; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4243 = 10'h3f6 == EXMEMALUOut[9:0] ? DMemory_1014 : _GEN_4242; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4244 = 10'h3f7 == EXMEMALUOut[9:0] ? DMemory_1015 : _GEN_4243; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4245 = 10'h3f8 == EXMEMALUOut[9:0] ? DMemory_1016 : _GEN_4244; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4246 = 10'h3f9 == EXMEMALUOut[9:0] ? DMemory_1017 : _GEN_4245; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4247 = 10'h3fa == EXMEMALUOut[9:0] ? DMemory_1018 : _GEN_4246; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4248 = 10'h3fb == EXMEMALUOut[9:0] ? DMemory_1019 : _GEN_4247; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4249 = 10'h3fc == EXMEMALUOut[9:0] ? DMemory_1020 : _GEN_4248; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4250 = 10'h3fd == EXMEMALUOut[9:0] ? DMemory_1021 : _GEN_4249; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4251 = 10'h3fe == EXMEMALUOut[9:0] ? DMemory_1022 : _GEN_4250; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4252 = 10'h3ff == EXMEMALUOut[9:0] ? DMemory_1023 : _GEN_4251; // @[CPU.scala 203:{18,18}]
  wire [31:0] _GEN_4253 = 10'h0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_0; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4254 = 10'h1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4255 = 10'h2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_2; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4256 = 10'h3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_3; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4257 = 10'h4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_4; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4258 = 10'h5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_5; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4259 = 10'h6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_6; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4260 = 10'h7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_7; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4261 = 10'h8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_8; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4262 = 10'h9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_9; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4263 = 10'ha == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_10; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4264 = 10'hb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_11; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4265 = 10'hc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_12; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4266 = 10'hd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_13; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4267 = 10'he == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_14; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4268 = 10'hf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_15; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4269 = 10'h10 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_16; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4270 = 10'h11 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_17; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4271 = 10'h12 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_18; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4272 = 10'h13 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_19; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4273 = 10'h14 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_20; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4274 = 10'h15 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_21; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4275 = 10'h16 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_22; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4276 = 10'h17 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_23; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4277 = 10'h18 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_24; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4278 = 10'h19 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_25; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4279 = 10'h1a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_26; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4280 = 10'h1b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_27; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4281 = 10'h1c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_28; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4282 = 10'h1d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_29; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4283 = 10'h1e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_30; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4284 = 10'h1f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_31; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4285 = 10'h20 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_32; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4286 = 10'h21 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_33; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4287 = 10'h22 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_34; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4288 = 10'h23 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_35; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4289 = 10'h24 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_36; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4290 = 10'h25 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_37; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4291 = 10'h26 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_38; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4292 = 10'h27 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_39; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4293 = 10'h28 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_40; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4294 = 10'h29 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_41; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4295 = 10'h2a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_42; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4296 = 10'h2b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_43; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4297 = 10'h2c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_44; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4298 = 10'h2d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_45; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4299 = 10'h2e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_46; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4300 = 10'h2f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_47; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4301 = 10'h30 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_48; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4302 = 10'h31 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_49; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4303 = 10'h32 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_50; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4304 = 10'h33 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_51; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4305 = 10'h34 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_52; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4306 = 10'h35 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_53; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4307 = 10'h36 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_54; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4308 = 10'h37 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_55; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4309 = 10'h38 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_56; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4310 = 10'h39 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_57; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4311 = 10'h3a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_58; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4312 = 10'h3b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_59; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4313 = 10'h3c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_60; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4314 = 10'h3d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_61; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4315 = 10'h3e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_62; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4316 = 10'h3f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_63; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4317 = 10'h40 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_64; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4318 = 10'h41 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_65; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4319 = 10'h42 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_66; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4320 = 10'h43 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_67; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4321 = 10'h44 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_68; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4322 = 10'h45 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_69; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4323 = 10'h46 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_70; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4324 = 10'h47 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_71; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4325 = 10'h48 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_72; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4326 = 10'h49 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_73; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4327 = 10'h4a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_74; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4328 = 10'h4b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_75; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4329 = 10'h4c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_76; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4330 = 10'h4d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_77; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4331 = 10'h4e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_78; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4332 = 10'h4f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_79; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4333 = 10'h50 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_80; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4334 = 10'h51 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_81; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4335 = 10'h52 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_82; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4336 = 10'h53 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_83; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4337 = 10'h54 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_84; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4338 = 10'h55 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_85; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4339 = 10'h56 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_86; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4340 = 10'h57 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_87; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4341 = 10'h58 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_88; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4342 = 10'h59 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_89; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4343 = 10'h5a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_90; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4344 = 10'h5b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_91; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4345 = 10'h5c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_92; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4346 = 10'h5d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_93; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4347 = 10'h5e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_94; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4348 = 10'h5f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_95; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4349 = 10'h60 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_96; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4350 = 10'h61 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_97; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4351 = 10'h62 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_98; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4352 = 10'h63 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_99; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4353 = 10'h64 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_100; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4354 = 10'h65 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_101; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4355 = 10'h66 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_102; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4356 = 10'h67 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_103; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4357 = 10'h68 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_104; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4358 = 10'h69 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_105; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4359 = 10'h6a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_106; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4360 = 10'h6b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_107; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4361 = 10'h6c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_108; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4362 = 10'h6d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_109; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4363 = 10'h6e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_110; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4364 = 10'h6f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_111; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4365 = 10'h70 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_112; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4366 = 10'h71 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_113; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4367 = 10'h72 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_114; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4368 = 10'h73 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_115; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4369 = 10'h74 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_116; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4370 = 10'h75 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_117; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4371 = 10'h76 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_118; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4372 = 10'h77 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_119; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4373 = 10'h78 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_120; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4374 = 10'h79 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_121; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4375 = 10'h7a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_122; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4376 = 10'h7b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_123; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4377 = 10'h7c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_124; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4378 = 10'h7d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_125; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4379 = 10'h7e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_126; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4380 = 10'h7f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_127; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4381 = 10'h80 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_128; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4382 = 10'h81 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_129; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4383 = 10'h82 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_130; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4384 = 10'h83 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_131; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4385 = 10'h84 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_132; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4386 = 10'h85 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_133; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4387 = 10'h86 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_134; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4388 = 10'h87 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_135; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4389 = 10'h88 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_136; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4390 = 10'h89 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_137; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4391 = 10'h8a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_138; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4392 = 10'h8b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_139; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4393 = 10'h8c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_140; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4394 = 10'h8d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_141; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4395 = 10'h8e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_142; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4396 = 10'h8f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_143; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4397 = 10'h90 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_144; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4398 = 10'h91 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_145; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4399 = 10'h92 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_146; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4400 = 10'h93 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_147; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4401 = 10'h94 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_148; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4402 = 10'h95 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_149; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4403 = 10'h96 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_150; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4404 = 10'h97 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_151; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4405 = 10'h98 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_152; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4406 = 10'h99 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_153; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4407 = 10'h9a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_154; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4408 = 10'h9b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_155; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4409 = 10'h9c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_156; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4410 = 10'h9d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_157; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4411 = 10'h9e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_158; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4412 = 10'h9f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_159; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4413 = 10'ha0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_160; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4414 = 10'ha1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_161; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4415 = 10'ha2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_162; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4416 = 10'ha3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_163; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4417 = 10'ha4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_164; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4418 = 10'ha5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_165; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4419 = 10'ha6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_166; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4420 = 10'ha7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_167; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4421 = 10'ha8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_168; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4422 = 10'ha9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_169; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4423 = 10'haa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_170; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4424 = 10'hab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_171; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4425 = 10'hac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_172; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4426 = 10'had == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_173; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4427 = 10'hae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_174; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4428 = 10'haf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_175; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4429 = 10'hb0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_176; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4430 = 10'hb1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_177; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4431 = 10'hb2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_178; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4432 = 10'hb3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_179; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4433 = 10'hb4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_180; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4434 = 10'hb5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_181; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4435 = 10'hb6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_182; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4436 = 10'hb7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_183; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4437 = 10'hb8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_184; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4438 = 10'hb9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_185; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4439 = 10'hba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_186; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4440 = 10'hbb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_187; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4441 = 10'hbc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_188; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4442 = 10'hbd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_189; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4443 = 10'hbe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_190; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4444 = 10'hbf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_191; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4445 = 10'hc0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_192; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4446 = 10'hc1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_193; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4447 = 10'hc2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_194; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4448 = 10'hc3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_195; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4449 = 10'hc4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_196; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4450 = 10'hc5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_197; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4451 = 10'hc6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_198; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4452 = 10'hc7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_199; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4453 = 10'hc8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_200; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4454 = 10'hc9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_201; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4455 = 10'hca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_202; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4456 = 10'hcb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_203; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4457 = 10'hcc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_204; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4458 = 10'hcd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_205; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4459 = 10'hce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_206; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4460 = 10'hcf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_207; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4461 = 10'hd0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_208; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4462 = 10'hd1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_209; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4463 = 10'hd2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_210; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4464 = 10'hd3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_211; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4465 = 10'hd4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_212; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4466 = 10'hd5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_213; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4467 = 10'hd6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_214; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4468 = 10'hd7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_215; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4469 = 10'hd8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_216; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4470 = 10'hd9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_217; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4471 = 10'hda == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_218; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4472 = 10'hdb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_219; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4473 = 10'hdc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_220; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4474 = 10'hdd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_221; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4475 = 10'hde == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_222; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4476 = 10'hdf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_223; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4477 = 10'he0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_224; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4478 = 10'he1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_225; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4479 = 10'he2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_226; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4480 = 10'he3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_227; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4481 = 10'he4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_228; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4482 = 10'he5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_229; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4483 = 10'he6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_230; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4484 = 10'he7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_231; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4485 = 10'he8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_232; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4486 = 10'he9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_233; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4487 = 10'hea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_234; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4488 = 10'heb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_235; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4489 = 10'hec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_236; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4490 = 10'hed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_237; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4491 = 10'hee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_238; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4492 = 10'hef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_239; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4493 = 10'hf0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_240; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4494 = 10'hf1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_241; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4495 = 10'hf2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_242; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4496 = 10'hf3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_243; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4497 = 10'hf4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_244; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4498 = 10'hf5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_245; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4499 = 10'hf6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_246; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4500 = 10'hf7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_247; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4501 = 10'hf8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_248; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4502 = 10'hf9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_249; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4503 = 10'hfa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_250; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4504 = 10'hfb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_251; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4505 = 10'hfc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_252; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4506 = 10'hfd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_253; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4507 = 10'hfe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_254; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4508 = 10'hff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_255; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4509 = 10'h100 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_256; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4510 = 10'h101 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_257; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4511 = 10'h102 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_258; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4512 = 10'h103 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_259; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4513 = 10'h104 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_260; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4514 = 10'h105 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_261; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4515 = 10'h106 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_262; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4516 = 10'h107 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_263; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4517 = 10'h108 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_264; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4518 = 10'h109 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_265; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4519 = 10'h10a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_266; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4520 = 10'h10b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_267; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4521 = 10'h10c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_268; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4522 = 10'h10d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_269; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4523 = 10'h10e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_270; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4524 = 10'h10f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_271; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4525 = 10'h110 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_272; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4526 = 10'h111 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_273; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4527 = 10'h112 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_274; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4528 = 10'h113 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_275; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4529 = 10'h114 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_276; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4530 = 10'h115 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_277; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4531 = 10'h116 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_278; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4532 = 10'h117 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_279; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4533 = 10'h118 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_280; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4534 = 10'h119 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_281; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4535 = 10'h11a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_282; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4536 = 10'h11b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_283; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4537 = 10'h11c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_284; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4538 = 10'h11d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_285; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4539 = 10'h11e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_286; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4540 = 10'h11f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_287; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4541 = 10'h120 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_288; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4542 = 10'h121 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_289; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4543 = 10'h122 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_290; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4544 = 10'h123 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_291; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4545 = 10'h124 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_292; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4546 = 10'h125 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_293; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4547 = 10'h126 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_294; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4548 = 10'h127 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_295; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4549 = 10'h128 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_296; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4550 = 10'h129 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_297; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4551 = 10'h12a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_298; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4552 = 10'h12b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_299; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4553 = 10'h12c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_300; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4554 = 10'h12d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_301; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4555 = 10'h12e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_302; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4556 = 10'h12f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_303; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4557 = 10'h130 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_304; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4558 = 10'h131 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_305; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4559 = 10'h132 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_306; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4560 = 10'h133 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_307; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4561 = 10'h134 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_308; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4562 = 10'h135 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_309; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4563 = 10'h136 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_310; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4564 = 10'h137 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_311; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4565 = 10'h138 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_312; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4566 = 10'h139 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_313; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4567 = 10'h13a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_314; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4568 = 10'h13b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_315; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4569 = 10'h13c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_316; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4570 = 10'h13d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_317; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4571 = 10'h13e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_318; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4572 = 10'h13f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_319; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4573 = 10'h140 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_320; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4574 = 10'h141 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_321; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4575 = 10'h142 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_322; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4576 = 10'h143 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_323; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4577 = 10'h144 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_324; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4578 = 10'h145 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_325; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4579 = 10'h146 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_326; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4580 = 10'h147 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_327; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4581 = 10'h148 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_328; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4582 = 10'h149 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_329; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4583 = 10'h14a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_330; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4584 = 10'h14b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_331; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4585 = 10'h14c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_332; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4586 = 10'h14d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_333; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4587 = 10'h14e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_334; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4588 = 10'h14f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_335; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4589 = 10'h150 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_336; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4590 = 10'h151 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_337; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4591 = 10'h152 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_338; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4592 = 10'h153 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_339; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4593 = 10'h154 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_340; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4594 = 10'h155 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_341; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4595 = 10'h156 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_342; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4596 = 10'h157 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_343; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4597 = 10'h158 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_344; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4598 = 10'h159 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_345; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4599 = 10'h15a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_346; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4600 = 10'h15b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_347; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4601 = 10'h15c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_348; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4602 = 10'h15d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_349; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4603 = 10'h15e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_350; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4604 = 10'h15f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_351; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4605 = 10'h160 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_352; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4606 = 10'h161 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_353; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4607 = 10'h162 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_354; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4608 = 10'h163 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_355; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4609 = 10'h164 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_356; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4610 = 10'h165 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_357; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4611 = 10'h166 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_358; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4612 = 10'h167 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_359; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4613 = 10'h168 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_360; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4614 = 10'h169 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_361; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4615 = 10'h16a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_362; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4616 = 10'h16b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_363; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4617 = 10'h16c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_364; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4618 = 10'h16d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_365; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4619 = 10'h16e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_366; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4620 = 10'h16f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_367; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4621 = 10'h170 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_368; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4622 = 10'h171 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_369; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4623 = 10'h172 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_370; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4624 = 10'h173 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_371; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4625 = 10'h174 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_372; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4626 = 10'h175 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_373; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4627 = 10'h176 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_374; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4628 = 10'h177 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_375; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4629 = 10'h178 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_376; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4630 = 10'h179 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_377; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4631 = 10'h17a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_378; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4632 = 10'h17b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_379; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4633 = 10'h17c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_380; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4634 = 10'h17d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_381; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4635 = 10'h17e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_382; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4636 = 10'h17f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_383; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4637 = 10'h180 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_384; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4638 = 10'h181 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_385; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4639 = 10'h182 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_386; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4640 = 10'h183 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_387; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4641 = 10'h184 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_388; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4642 = 10'h185 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_389; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4643 = 10'h186 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_390; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4644 = 10'h187 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_391; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4645 = 10'h188 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_392; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4646 = 10'h189 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_393; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4647 = 10'h18a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_394; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4648 = 10'h18b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_395; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4649 = 10'h18c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_396; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4650 = 10'h18d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_397; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4651 = 10'h18e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_398; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4652 = 10'h18f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_399; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4653 = 10'h190 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_400; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4654 = 10'h191 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_401; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4655 = 10'h192 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_402; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4656 = 10'h193 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_403; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4657 = 10'h194 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_404; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4658 = 10'h195 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_405; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4659 = 10'h196 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_406; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4660 = 10'h197 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_407; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4661 = 10'h198 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_408; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4662 = 10'h199 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_409; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4663 = 10'h19a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_410; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4664 = 10'h19b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_411; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4665 = 10'h19c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_412; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4666 = 10'h19d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_413; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4667 = 10'h19e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_414; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4668 = 10'h19f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_415; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4669 = 10'h1a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_416; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4670 = 10'h1a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_417; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4671 = 10'h1a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_418; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4672 = 10'h1a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_419; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4673 = 10'h1a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_420; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4674 = 10'h1a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_421; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4675 = 10'h1a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_422; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4676 = 10'h1a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_423; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4677 = 10'h1a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_424; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4678 = 10'h1a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_425; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4679 = 10'h1aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_426; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4680 = 10'h1ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_427; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4681 = 10'h1ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_428; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4682 = 10'h1ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_429; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4683 = 10'h1ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_430; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4684 = 10'h1af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_431; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4685 = 10'h1b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_432; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4686 = 10'h1b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_433; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4687 = 10'h1b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_434; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4688 = 10'h1b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_435; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4689 = 10'h1b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_436; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4690 = 10'h1b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_437; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4691 = 10'h1b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_438; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4692 = 10'h1b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_439; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4693 = 10'h1b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_440; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4694 = 10'h1b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_441; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4695 = 10'h1ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_442; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4696 = 10'h1bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_443; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4697 = 10'h1bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_444; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4698 = 10'h1bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_445; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4699 = 10'h1be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_446; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4700 = 10'h1bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_447; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4701 = 10'h1c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_448; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4702 = 10'h1c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_449; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4703 = 10'h1c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_450; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4704 = 10'h1c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_451; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4705 = 10'h1c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_452; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4706 = 10'h1c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_453; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4707 = 10'h1c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_454; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4708 = 10'h1c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_455; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4709 = 10'h1c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_456; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4710 = 10'h1c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_457; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4711 = 10'h1ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_458; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4712 = 10'h1cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_459; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4713 = 10'h1cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_460; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4714 = 10'h1cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_461; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4715 = 10'h1ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_462; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4716 = 10'h1cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_463; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4717 = 10'h1d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_464; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4718 = 10'h1d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_465; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4719 = 10'h1d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_466; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4720 = 10'h1d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_467; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4721 = 10'h1d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_468; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4722 = 10'h1d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_469; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4723 = 10'h1d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_470; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4724 = 10'h1d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_471; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4725 = 10'h1d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_472; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4726 = 10'h1d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_473; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4727 = 10'h1da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_474; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4728 = 10'h1db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_475; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4729 = 10'h1dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_476; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4730 = 10'h1dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_477; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4731 = 10'h1de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_478; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4732 = 10'h1df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_479; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4733 = 10'h1e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_480; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4734 = 10'h1e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_481; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4735 = 10'h1e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_482; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4736 = 10'h1e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_483; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4737 = 10'h1e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_484; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4738 = 10'h1e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_485; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4739 = 10'h1e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_486; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4740 = 10'h1e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_487; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4741 = 10'h1e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_488; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4742 = 10'h1e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_489; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4743 = 10'h1ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_490; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4744 = 10'h1eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_491; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4745 = 10'h1ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_492; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4746 = 10'h1ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_493; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4747 = 10'h1ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_494; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4748 = 10'h1ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_495; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4749 = 10'h1f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_496; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4750 = 10'h1f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_497; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4751 = 10'h1f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_498; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4752 = 10'h1f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_499; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4753 = 10'h1f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_500; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4754 = 10'h1f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_501; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4755 = 10'h1f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_502; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4756 = 10'h1f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_503; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4757 = 10'h1f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_504; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4758 = 10'h1f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_505; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4759 = 10'h1fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_506; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4760 = 10'h1fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_507; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4761 = 10'h1fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_508; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4762 = 10'h1fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_509; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4763 = 10'h1fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_510; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4764 = 10'h1ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_511; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4765 = 10'h200 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_512; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4766 = 10'h201 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_513; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4767 = 10'h202 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_514; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4768 = 10'h203 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_515; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4769 = 10'h204 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_516; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4770 = 10'h205 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_517; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4771 = 10'h206 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_518; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4772 = 10'h207 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_519; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4773 = 10'h208 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_520; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4774 = 10'h209 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_521; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4775 = 10'h20a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_522; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4776 = 10'h20b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_523; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4777 = 10'h20c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_524; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4778 = 10'h20d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_525; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4779 = 10'h20e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_526; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4780 = 10'h20f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_527; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4781 = 10'h210 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_528; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4782 = 10'h211 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_529; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4783 = 10'h212 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_530; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4784 = 10'h213 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_531; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4785 = 10'h214 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_532; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4786 = 10'h215 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_533; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4787 = 10'h216 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_534; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4788 = 10'h217 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_535; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4789 = 10'h218 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_536; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4790 = 10'h219 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_537; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4791 = 10'h21a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_538; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4792 = 10'h21b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_539; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4793 = 10'h21c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_540; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4794 = 10'h21d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_541; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4795 = 10'h21e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_542; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4796 = 10'h21f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_543; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4797 = 10'h220 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_544; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4798 = 10'h221 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_545; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4799 = 10'h222 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_546; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4800 = 10'h223 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_547; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4801 = 10'h224 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_548; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4802 = 10'h225 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_549; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4803 = 10'h226 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_550; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4804 = 10'h227 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_551; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4805 = 10'h228 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_552; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4806 = 10'h229 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_553; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4807 = 10'h22a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_554; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4808 = 10'h22b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_555; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4809 = 10'h22c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_556; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4810 = 10'h22d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_557; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4811 = 10'h22e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_558; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4812 = 10'h22f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_559; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4813 = 10'h230 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_560; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4814 = 10'h231 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_561; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4815 = 10'h232 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_562; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4816 = 10'h233 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_563; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4817 = 10'h234 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_564; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4818 = 10'h235 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_565; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4819 = 10'h236 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_566; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4820 = 10'h237 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_567; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4821 = 10'h238 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_568; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4822 = 10'h239 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_569; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4823 = 10'h23a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_570; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4824 = 10'h23b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_571; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4825 = 10'h23c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_572; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4826 = 10'h23d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_573; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4827 = 10'h23e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_574; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4828 = 10'h23f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_575; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4829 = 10'h240 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_576; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4830 = 10'h241 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_577; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4831 = 10'h242 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_578; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4832 = 10'h243 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_579; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4833 = 10'h244 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_580; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4834 = 10'h245 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_581; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4835 = 10'h246 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_582; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4836 = 10'h247 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_583; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4837 = 10'h248 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_584; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4838 = 10'h249 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_585; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4839 = 10'h24a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_586; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4840 = 10'h24b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_587; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4841 = 10'h24c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_588; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4842 = 10'h24d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_589; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4843 = 10'h24e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_590; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4844 = 10'h24f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_591; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4845 = 10'h250 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_592; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4846 = 10'h251 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_593; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4847 = 10'h252 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_594; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4848 = 10'h253 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_595; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4849 = 10'h254 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_596; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4850 = 10'h255 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_597; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4851 = 10'h256 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_598; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4852 = 10'h257 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_599; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4853 = 10'h258 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_600; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4854 = 10'h259 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_601; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4855 = 10'h25a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_602; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4856 = 10'h25b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_603; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4857 = 10'h25c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_604; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4858 = 10'h25d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_605; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4859 = 10'h25e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_606; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4860 = 10'h25f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_607; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4861 = 10'h260 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_608; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4862 = 10'h261 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_609; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4863 = 10'h262 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_610; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4864 = 10'h263 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_611; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4865 = 10'h264 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_612; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4866 = 10'h265 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_613; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4867 = 10'h266 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_614; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4868 = 10'h267 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_615; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4869 = 10'h268 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_616; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4870 = 10'h269 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_617; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4871 = 10'h26a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_618; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4872 = 10'h26b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_619; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4873 = 10'h26c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_620; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4874 = 10'h26d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_621; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4875 = 10'h26e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_622; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4876 = 10'h26f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_623; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4877 = 10'h270 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_624; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4878 = 10'h271 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_625; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4879 = 10'h272 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_626; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4880 = 10'h273 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_627; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4881 = 10'h274 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_628; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4882 = 10'h275 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_629; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4883 = 10'h276 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_630; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4884 = 10'h277 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_631; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4885 = 10'h278 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_632; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4886 = 10'h279 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_633; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4887 = 10'h27a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_634; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4888 = 10'h27b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_635; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4889 = 10'h27c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_636; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4890 = 10'h27d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_637; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4891 = 10'h27e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_638; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4892 = 10'h27f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_639; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4893 = 10'h280 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_640; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4894 = 10'h281 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_641; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4895 = 10'h282 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_642; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4896 = 10'h283 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_643; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4897 = 10'h284 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_644; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4898 = 10'h285 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_645; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4899 = 10'h286 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_646; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4900 = 10'h287 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_647; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4901 = 10'h288 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_648; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4902 = 10'h289 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_649; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4903 = 10'h28a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_650; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4904 = 10'h28b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_651; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4905 = 10'h28c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_652; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4906 = 10'h28d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_653; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4907 = 10'h28e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_654; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4908 = 10'h28f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_655; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4909 = 10'h290 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_656; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4910 = 10'h291 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_657; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4911 = 10'h292 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_658; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4912 = 10'h293 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_659; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4913 = 10'h294 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_660; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4914 = 10'h295 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_661; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4915 = 10'h296 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_662; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4916 = 10'h297 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_663; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4917 = 10'h298 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_664; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4918 = 10'h299 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_665; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4919 = 10'h29a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_666; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4920 = 10'h29b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_667; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4921 = 10'h29c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_668; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4922 = 10'h29d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_669; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4923 = 10'h29e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_670; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4924 = 10'h29f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_671; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4925 = 10'h2a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_672; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4926 = 10'h2a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_673; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4927 = 10'h2a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_674; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4928 = 10'h2a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_675; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4929 = 10'h2a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_676; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4930 = 10'h2a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_677; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4931 = 10'h2a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_678; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4932 = 10'h2a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_679; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4933 = 10'h2a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_680; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4934 = 10'h2a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_681; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4935 = 10'h2aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_682; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4936 = 10'h2ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_683; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4937 = 10'h2ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_684; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4938 = 10'h2ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_685; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4939 = 10'h2ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_686; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4940 = 10'h2af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_687; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4941 = 10'h2b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_688; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4942 = 10'h2b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_689; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4943 = 10'h2b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_690; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4944 = 10'h2b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_691; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4945 = 10'h2b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_692; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4946 = 10'h2b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_693; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4947 = 10'h2b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_694; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4948 = 10'h2b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_695; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4949 = 10'h2b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_696; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4950 = 10'h2b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_697; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4951 = 10'h2ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_698; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4952 = 10'h2bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_699; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4953 = 10'h2bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_700; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4954 = 10'h2bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_701; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4955 = 10'h2be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_702; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4956 = 10'h2bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_703; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4957 = 10'h2c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_704; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4958 = 10'h2c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_705; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4959 = 10'h2c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_706; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4960 = 10'h2c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_707; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4961 = 10'h2c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_708; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4962 = 10'h2c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_709; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4963 = 10'h2c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_710; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4964 = 10'h2c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_711; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4965 = 10'h2c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_712; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4966 = 10'h2c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_713; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4967 = 10'h2ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_714; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4968 = 10'h2cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_715; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4969 = 10'h2cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_716; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4970 = 10'h2cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_717; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4971 = 10'h2ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_718; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4972 = 10'h2cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_719; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4973 = 10'h2d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_720; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4974 = 10'h2d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_721; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4975 = 10'h2d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_722; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4976 = 10'h2d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_723; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4977 = 10'h2d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_724; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4978 = 10'h2d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_725; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4979 = 10'h2d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_726; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4980 = 10'h2d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_727; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4981 = 10'h2d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_728; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4982 = 10'h2d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_729; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4983 = 10'h2da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_730; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4984 = 10'h2db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_731; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4985 = 10'h2dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_732; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4986 = 10'h2dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_733; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4987 = 10'h2de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_734; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4988 = 10'h2df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_735; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4989 = 10'h2e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_736; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4990 = 10'h2e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_737; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4991 = 10'h2e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_738; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4992 = 10'h2e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_739; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4993 = 10'h2e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_740; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4994 = 10'h2e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_741; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4995 = 10'h2e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_742; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4996 = 10'h2e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_743; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4997 = 10'h2e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_744; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4998 = 10'h2e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_745; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_4999 = 10'h2ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_746; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5000 = 10'h2eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_747; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5001 = 10'h2ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_748; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5002 = 10'h2ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_749; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5003 = 10'h2ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_750; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5004 = 10'h2ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_751; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5005 = 10'h2f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_752; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5006 = 10'h2f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_753; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5007 = 10'h2f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_754; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5008 = 10'h2f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_755; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5009 = 10'h2f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_756; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5010 = 10'h2f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_757; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5011 = 10'h2f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_758; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5012 = 10'h2f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_759; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5013 = 10'h2f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_760; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5014 = 10'h2f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_761; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5015 = 10'h2fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_762; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5016 = 10'h2fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_763; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5017 = 10'h2fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_764; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5018 = 10'h2fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_765; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5019 = 10'h2fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_766; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5020 = 10'h2ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_767; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5021 = 10'h300 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_768; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5022 = 10'h301 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_769; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5023 = 10'h302 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_770; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5024 = 10'h303 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_771; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5025 = 10'h304 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_772; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5026 = 10'h305 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_773; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5027 = 10'h306 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_774; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5028 = 10'h307 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_775; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5029 = 10'h308 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_776; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5030 = 10'h309 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_777; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5031 = 10'h30a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_778; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5032 = 10'h30b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_779; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5033 = 10'h30c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_780; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5034 = 10'h30d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_781; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5035 = 10'h30e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_782; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5036 = 10'h30f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_783; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5037 = 10'h310 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_784; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5038 = 10'h311 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_785; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5039 = 10'h312 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_786; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5040 = 10'h313 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_787; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5041 = 10'h314 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_788; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5042 = 10'h315 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_789; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5043 = 10'h316 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_790; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5044 = 10'h317 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_791; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5045 = 10'h318 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_792; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5046 = 10'h319 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_793; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5047 = 10'h31a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_794; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5048 = 10'h31b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_795; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5049 = 10'h31c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_796; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5050 = 10'h31d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_797; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5051 = 10'h31e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_798; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5052 = 10'h31f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_799; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5053 = 10'h320 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_800; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5054 = 10'h321 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_801; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5055 = 10'h322 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_802; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5056 = 10'h323 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_803; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5057 = 10'h324 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_804; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5058 = 10'h325 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_805; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5059 = 10'h326 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_806; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5060 = 10'h327 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_807; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5061 = 10'h328 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_808; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5062 = 10'h329 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_809; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5063 = 10'h32a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_810; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5064 = 10'h32b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_811; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5065 = 10'h32c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_812; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5066 = 10'h32d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_813; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5067 = 10'h32e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_814; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5068 = 10'h32f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_815; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5069 = 10'h330 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_816; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5070 = 10'h331 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_817; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5071 = 10'h332 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_818; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5072 = 10'h333 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_819; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5073 = 10'h334 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_820; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5074 = 10'h335 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_821; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5075 = 10'h336 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_822; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5076 = 10'h337 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_823; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5077 = 10'h338 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_824; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5078 = 10'h339 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_825; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5079 = 10'h33a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_826; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5080 = 10'h33b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_827; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5081 = 10'h33c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_828; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5082 = 10'h33d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_829; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5083 = 10'h33e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_830; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5084 = 10'h33f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_831; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5085 = 10'h340 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_832; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5086 = 10'h341 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_833; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5087 = 10'h342 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_834; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5088 = 10'h343 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_835; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5089 = 10'h344 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_836; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5090 = 10'h345 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_837; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5091 = 10'h346 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_838; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5092 = 10'h347 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_839; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5093 = 10'h348 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_840; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5094 = 10'h349 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_841; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5095 = 10'h34a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_842; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5096 = 10'h34b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_843; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5097 = 10'h34c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_844; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5098 = 10'h34d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_845; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5099 = 10'h34e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_846; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5100 = 10'h34f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_847; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5101 = 10'h350 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_848; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5102 = 10'h351 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_849; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5103 = 10'h352 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_850; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5104 = 10'h353 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_851; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5105 = 10'h354 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_852; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5106 = 10'h355 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_853; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5107 = 10'h356 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_854; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5108 = 10'h357 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_855; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5109 = 10'h358 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_856; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5110 = 10'h359 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_857; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5111 = 10'h35a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_858; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5112 = 10'h35b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_859; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5113 = 10'h35c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_860; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5114 = 10'h35d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_861; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5115 = 10'h35e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_862; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5116 = 10'h35f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_863; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5117 = 10'h360 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_864; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5118 = 10'h361 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_865; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5119 = 10'h362 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_866; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5120 = 10'h363 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_867; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5121 = 10'h364 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_868; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5122 = 10'h365 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_869; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5123 = 10'h366 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_870; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5124 = 10'h367 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_871; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5125 = 10'h368 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_872; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5126 = 10'h369 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_873; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5127 = 10'h36a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_874; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5128 = 10'h36b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_875; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5129 = 10'h36c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_876; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5130 = 10'h36d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_877; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5131 = 10'h36e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_878; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5132 = 10'h36f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_879; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5133 = 10'h370 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_880; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5134 = 10'h371 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_881; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5135 = 10'h372 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_882; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5136 = 10'h373 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_883; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5137 = 10'h374 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_884; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5138 = 10'h375 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_885; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5139 = 10'h376 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_886; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5140 = 10'h377 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_887; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5141 = 10'h378 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_888; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5142 = 10'h379 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_889; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5143 = 10'h37a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_890; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5144 = 10'h37b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_891; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5145 = 10'h37c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_892; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5146 = 10'h37d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_893; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5147 = 10'h37e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_894; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5148 = 10'h37f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_895; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5149 = 10'h380 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_896; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5150 = 10'h381 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_897; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5151 = 10'h382 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_898; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5152 = 10'h383 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_899; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5153 = 10'h384 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_900; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5154 = 10'h385 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_901; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5155 = 10'h386 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_902; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5156 = 10'h387 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_903; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5157 = 10'h388 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_904; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5158 = 10'h389 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_905; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5159 = 10'h38a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_906; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5160 = 10'h38b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_907; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5161 = 10'h38c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_908; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5162 = 10'h38d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_909; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5163 = 10'h38e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_910; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5164 = 10'h38f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_911; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5165 = 10'h390 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_912; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5166 = 10'h391 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_913; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5167 = 10'h392 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_914; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5168 = 10'h393 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_915; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5169 = 10'h394 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_916; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5170 = 10'h395 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_917; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5171 = 10'h396 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_918; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5172 = 10'h397 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_919; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5173 = 10'h398 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_920; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5174 = 10'h399 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_921; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5175 = 10'h39a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_922; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5176 = 10'h39b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_923; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5177 = 10'h39c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_924; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5178 = 10'h39d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_925; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5179 = 10'h39e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_926; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5180 = 10'h39f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_927; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5181 = 10'h3a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_928; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5182 = 10'h3a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_929; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5183 = 10'h3a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_930; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5184 = 10'h3a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_931; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5185 = 10'h3a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_932; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5186 = 10'h3a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_933; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5187 = 10'h3a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_934; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5188 = 10'h3a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_935; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5189 = 10'h3a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_936; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5190 = 10'h3a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_937; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5191 = 10'h3aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_938; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5192 = 10'h3ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_939; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5193 = 10'h3ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_940; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5194 = 10'h3ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_941; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5195 = 10'h3ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_942; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5196 = 10'h3af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_943; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5197 = 10'h3b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_944; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5198 = 10'h3b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_945; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5199 = 10'h3b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_946; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5200 = 10'h3b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_947; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5201 = 10'h3b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_948; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5202 = 10'h3b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_949; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5203 = 10'h3b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_950; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5204 = 10'h3b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_951; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5205 = 10'h3b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_952; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5206 = 10'h3b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_953; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5207 = 10'h3ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_954; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5208 = 10'h3bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_955; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5209 = 10'h3bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_956; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5210 = 10'h3bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_957; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5211 = 10'h3be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_958; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5212 = 10'h3bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_959; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5213 = 10'h3c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_960; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5214 = 10'h3c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_961; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5215 = 10'h3c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_962; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5216 = 10'h3c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_963; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5217 = 10'h3c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_964; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5218 = 10'h3c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_965; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5219 = 10'h3c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_966; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5220 = 10'h3c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_967; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5221 = 10'h3c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_968; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5222 = 10'h3c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_969; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5223 = 10'h3ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_970; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5224 = 10'h3cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_971; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5225 = 10'h3cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_972; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5226 = 10'h3cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_973; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5227 = 10'h3ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_974; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5228 = 10'h3cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_975; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5229 = 10'h3d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_976; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5230 = 10'h3d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_977; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5231 = 10'h3d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_978; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5232 = 10'h3d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_979; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5233 = 10'h3d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_980; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5234 = 10'h3d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_981; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5235 = 10'h3d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_982; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5236 = 10'h3d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_983; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5237 = 10'h3d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_984; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5238 = 10'h3d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_985; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5239 = 10'h3da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_986; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5240 = 10'h3db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_987; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5241 = 10'h3dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_988; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5242 = 10'h3dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_989; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5243 = 10'h3de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_990; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5244 = 10'h3df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_991; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5245 = 10'h3e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_992; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5246 = 10'h3e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_993; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5247 = 10'h3e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_994; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5248 = 10'h3e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_995; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5249 = 10'h3e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_996; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5250 = 10'h3e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_997; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5251 = 10'h3e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_998; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5252 = 10'h3e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_999; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5253 = 10'h3e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1000; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5254 = 10'h3e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1001; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5255 = 10'h3ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1002; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5256 = 10'h3eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1003; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5257 = 10'h3ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1004; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5258 = 10'h3ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1005; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5259 = 10'h3ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1006; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5260 = 10'h3ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1007; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5261 = 10'h3f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1008; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5262 = 10'h3f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1009; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5263 = 10'h3f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1010; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5264 = 10'h3f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1011; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5265 = 10'h3f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1012; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5266 = 10'h3f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1013; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5267 = 10'h3f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1014; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5268 = 10'h3f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1015; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5269 = 10'h3f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1016; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5270 = 10'h3f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1017; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5271 = 10'h3fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1018; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5272 = 10'h3fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1019; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5273 = 10'h3fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1020; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5274 = 10'h3fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1021; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5275 = 10'h3fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1022; // @[CPU.scala 205:{37,37} 52:20]
  wire [31:0] _GEN_5276 = 10'h3ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1023; // @[CPU.scala 205:{37,37} 52:20]
  assign io_rvfi_valid = 1'h0; // @[CPU.scala 223:17]
  assign io_rvfi_insn = MEMWBIR; // @[CPU.scala 222:16]
  assign io_rvfi_pc_rdata = CurPC; // @[CPU.scala 226:20]
  assign io_rvfi_pc_wdata = PC; // @[CPU.scala 228:20]
  assign io_rvfi_rs1_addr = io_rvfi_rst ? IFIDIR[19:15] : IFIDIR[19:15]; // @[CPU.scala 61:21 64:13 81:13]
  assign io_rvfi_rs2_addr = io_rvfi_rst ? IFIDIR[24:20] : IFIDIR[24:20]; // @[CPU.scala 61:21 65:13 82:13]
  assign io_rvfi_rs1_rdata = IDEXA; // @[CPU.scala 234:21]
  assign io_rvfi_rs2_rdata = IDEXB; // @[CPU.scala 236:21]
  assign io_rvfi_rd_addr = io_rvfi_rst ? MEMWBIR[11:7] : MEMWBIR[11:7]; // @[CPU.scala 61:21 70:13 87:13]
  assign io_rvfi_rd_wdata = MEMWBValue; // @[CPU.scala 219:20]
  assign io_rvfi_mem_addr = EXMEMALUOut[31:0]; // @[CPU.scala 240:20]
  assign io_rvfi_mem_rdata = MEMWBValue; // @[CPU.scala 242:21]
  assign io_rvfi_mem_wdata = {{32'd0}, DMemory_1}; // @[CPU.scala 244:21]
  assign io_rvfi_regs_0 = Regs_0; // @[CPU.scala 221:16]
  assign io_rvfi_regs_1 = Regs_1; // @[CPU.scala 221:16]
  assign io_rvfi_regs_2 = Regs_2; // @[CPU.scala 221:16]
  assign io_rvfi_regs_3 = Regs_3; // @[CPU.scala 221:16]
  assign io_rvfi_regs_4 = Regs_4; // @[CPU.scala 221:16]
  assign io_rvfi_regs_5 = Regs_5; // @[CPU.scala 221:16]
  assign io_rvfi_regs_6 = Regs_6; // @[CPU.scala 221:16]
  assign io_rvfi_regs_7 = Regs_7; // @[CPU.scala 221:16]
  assign io_rvfi_regs_8 = Regs_8; // @[CPU.scala 221:16]
  assign io_rvfi_regs_9 = Regs_9; // @[CPU.scala 221:16]
  assign io_rvfi_regs_10 = Regs_10; // @[CPU.scala 221:16]
  assign io_rvfi_regs_11 = Regs_11; // @[CPU.scala 221:16]
  assign io_rvfi_regs_12 = Regs_12; // @[CPU.scala 221:16]
  assign io_rvfi_regs_13 = Regs_13; // @[CPU.scala 221:16]
  assign io_rvfi_regs_14 = Regs_14; // @[CPU.scala 221:16]
  assign io_rvfi_regs_15 = Regs_15; // @[CPU.scala 221:16]
  assign io_rvfi_regs_16 = Regs_16; // @[CPU.scala 221:16]
  assign io_rvfi_regs_17 = Regs_17; // @[CPU.scala 221:16]
  assign io_rvfi_regs_18 = Regs_18; // @[CPU.scala 221:16]
  assign io_rvfi_regs_19 = Regs_19; // @[CPU.scala 221:16]
  assign io_rvfi_regs_20 = Regs_20; // @[CPU.scala 221:16]
  assign io_rvfi_regs_21 = Regs_21; // @[CPU.scala 221:16]
  assign io_rvfi_regs_22 = Regs_22; // @[CPU.scala 221:16]
  assign io_rvfi_regs_23 = Regs_23; // @[CPU.scala 221:16]
  assign io_rvfi_regs_24 = Regs_24; // @[CPU.scala 221:16]
  assign io_rvfi_regs_25 = Regs_25; // @[CPU.scala 221:16]
  assign io_rvfi_regs_26 = Regs_26; // @[CPU.scala 221:16]
  assign io_rvfi_regs_27 = Regs_27; // @[CPU.scala 221:16]
  assign io_rvfi_regs_28 = Regs_28; // @[CPU.scala 221:16]
  assign io_rvfi_regs_29 = Regs_29; // @[CPU.scala 221:16]
  assign io_rvfi_regs_30 = Regs_30; // @[CPU.scala 221:16]
  assign io_rvfi_regs_31 = Regs_31; // @[CPU.scala 221:16]
  always @(posedge clock) begin
    if (reset) begin // @[CPU.scala 48:19]
      PC <= 64'h0; // @[CPU.scala 48:19]
    end else if (!(io_rvfi_rst)) begin // @[CPU.scala 61:21]
      if (~stall) begin // @[CPU.scala 121:27]
        if (~takeBranch) begin // @[CPU.scala 122:34]
          PC <= _PC_T_1; // @[CPU.scala 126:12]
        end else begin
          PC <= branchTarget; // @[CPU.scala 142:12]
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h0 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_0 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h0 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_0 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h0 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_0 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h1 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_1 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h1 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_1 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h1 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_1 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h2 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_2 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h2 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_2 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h2 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_2 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h3 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_3 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h3 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_3 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h3 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_3 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h4 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_4 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h4 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_4 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h4 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_4 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h5 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_5 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h5 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_5 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h5 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_5 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h6 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_6 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h6 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_6 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h6 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_6 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h7 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_7 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h7 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_7 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h7 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_7 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h8 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_8 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h8 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_8 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h8 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_8 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h9 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_9 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h9 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_9 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h9 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_9 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'ha == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_10 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'ha == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_10 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'ha == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_10 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'hb == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_11 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'hb == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_11 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'hb == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_11 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'hc == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_12 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'hc == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_12 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'hc == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_12 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'hd == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_13 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'hd == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_13 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'hd == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_13 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'he == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_14 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'he == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_14 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'he == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_14 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'hf == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_15 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'hf == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_15 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'hf == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_15 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h10 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_16 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h10 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_16 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h10 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_16 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h11 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_17 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h11 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_17 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h11 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_17 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h12 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_18 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h12 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_18 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h12 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_18 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h13 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_19 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h13 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_19 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h13 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_19 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h14 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_20 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h14 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_20 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h14 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_20 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h15 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_21 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h15 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_21 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h15 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_21 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h16 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_22 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h16 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_22 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h16 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_22 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h17 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_23 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h17 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_23 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h17 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_23 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h18 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_24 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h18 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_24 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h18 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_24 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h19 == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_25 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h19 == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_25 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h19 == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_25 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h1a == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_26 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h1a == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_26 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h1a == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_26 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h1b == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_27 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h1b == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_27 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h1b == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_27 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h1c == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_28 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h1c == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_28 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h1c == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_28 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h1d == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_29 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h1d == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_29 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h1d == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_29 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h1e == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_30 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h1e == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_30 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h1e == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_30 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (5'h1f == io_rvfi_rs2_addr_in) begin // @[CPU.scala 63:31]
        Regs_31 <= io_rvfi_rs2_rdata_in; // @[CPU.scala 63:31]
      end else if (5'h1f == io_rvfi_rs1_addr_in) begin // @[CPU.scala 62:31]
        Regs_31 <= io_rvfi_rs1_rdata_in; // @[CPU.scala 62:31]
      end
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[CPU.scala 214:74]
      if (5'h1f == MEMWBrd) begin // @[CPU.scala 215:21]
        Regs_31 <= MEMWBValue; // @[CPU.scala 215:21]
      end
    end
    if (!(io_rvfi_rst)) begin // @[CPU.scala 61:21]
      if (~stall) begin // @[CPU.scala 121:27]
        if (bypassAFromEX) begin // @[CPU.scala 148:27]
          IDEXA <= _A_T_1; // @[CPU.scala 150:11]
        end else if (bypassAFromMEM) begin // @[CPU.scala 151:34]
          IDEXA <= EXMEMALUOut; // @[CPU.scala 153:11]
        end else begin
          IDEXA <= _GEN_3173;
        end
      end else begin
        IDEXA <= 64'h0;
      end
    end
    if (!(io_rvfi_rst)) begin // @[CPU.scala 61:21]
      if (~stall) begin // @[CPU.scala 121:27]
        if (bypassBFromEX) begin // @[CPU.scala 161:27]
          IDEXB <= _B_T_1; // @[CPU.scala 163:11]
        end else if (bypassBFromMEM) begin // @[CPU.scala 164:34]
          IDEXB <= EXMEMALUOut; // @[CPU.scala 166:11]
        end else begin
          IDEXB <= _GEN_3211;
        end
      end else begin
        IDEXB <= 64'h0;
      end
    end
    if (!(io_rvfi_rst)) begin // @[CPU.scala 61:21]
      EXMEMB <= IDEXB; // @[CPU.scala 197:12]
    end
    if (!(io_rvfi_rst)) begin // @[CPU.scala 61:21]
      if (_stall_T_9) begin // @[CPU.scala 182:25]
        EXMEMALUOut <= _EXMEMALUOut_T_6; // @[CPU.scala 183:19]
      end else if (IDEXop == 7'h23) begin // @[CPU.scala 184:31]
        EXMEMALUOut <= _EXMEMALUOut_T_15; // @[CPU.scala 185:19]
      end else if (_bypassAFromEX_T_3) begin // @[CPU.scala 189:34]
        EXMEMALUOut <= _A_T_1; // @[CPU.scala 192:19]
      end
    end
    if (!(io_rvfi_rst)) begin // @[CPU.scala 61:21]
      if (_bypassAFromMEM_T_3) begin // @[CPU.scala 200:29]
        MEMWBValue <= EXMEMALUOut; // @[CPU.scala 201:18]
      end else if (_stall_T) begin // @[CPU.scala 202:32]
        MEMWBValue <= {{32'd0}, _GEN_4252}; // @[CPU.scala 203:18]
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_0 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_0 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_0 <= _GEN_4253;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1 <= _GEN_4254;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_2 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_2 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_2 <= _GEN_4255;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_3 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_3 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_3 <= _GEN_4256;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_4 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_4 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_4 <= _GEN_4257;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_5 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_5 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_5 <= _GEN_4258;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_6 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_6 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_6 <= _GEN_4259;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_7 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_7 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_7 <= _GEN_4260;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_8 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_8 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_8 <= _GEN_4261;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_9 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_9 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_9 <= _GEN_4262;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'ha == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_10 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'ha == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_10 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_10 <= _GEN_4263;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_11 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_11 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_11 <= _GEN_4264;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_12 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_12 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_12 <= _GEN_4265;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_13 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_13 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_13 <= _GEN_4266;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'he == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_14 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'he == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_14 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_14 <= _GEN_4267;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hf == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_15 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hf == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_15 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_15 <= _GEN_4268;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h10 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_16 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h10 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_16 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_16 <= _GEN_4269;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h11 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_17 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h11 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_17 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_17 <= _GEN_4270;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h12 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_18 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h12 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_18 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_18 <= _GEN_4271;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h13 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_19 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h13 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_19 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_19 <= _GEN_4272;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h14 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_20 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h14 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_20 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_20 <= _GEN_4273;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h15 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_21 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h15 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_21 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_21 <= _GEN_4274;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h16 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_22 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h16 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_22 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_22 <= _GEN_4275;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h17 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_23 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h17 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_23 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_23 <= _GEN_4276;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h18 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_24 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h18 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_24 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_24 <= _GEN_4277;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h19 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_25 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h19 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_25 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_25 <= _GEN_4278;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_26 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_26 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_26 <= _GEN_4279;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_27 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_27 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_27 <= _GEN_4280;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_28 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_28 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_28 <= _GEN_4281;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_29 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_29 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_29 <= _GEN_4282;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_30 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_30 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_30 <= _GEN_4283;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_31 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_31 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_31 <= _GEN_4284;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h20 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_32 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h20 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_32 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_32 <= _GEN_4285;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h21 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_33 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h21 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_33 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_33 <= _GEN_4286;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h22 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_34 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h22 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_34 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_34 <= _GEN_4287;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h23 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_35 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h23 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_35 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_35 <= _GEN_4288;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h24 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_36 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h24 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_36 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_36 <= _GEN_4289;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h25 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_37 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h25 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_37 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_37 <= _GEN_4290;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h26 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_38 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h26 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_38 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_38 <= _GEN_4291;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h27 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_39 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h27 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_39 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_39 <= _GEN_4292;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h28 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_40 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h28 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_40 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_40 <= _GEN_4293;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h29 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_41 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h29 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_41 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_41 <= _GEN_4294;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_42 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_42 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_42 <= _GEN_4295;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_43 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_43 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_43 <= _GEN_4296;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_44 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_44 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_44 <= _GEN_4297;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_45 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_45 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_45 <= _GEN_4298;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_46 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_46 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_46 <= _GEN_4299;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_47 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_47 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_47 <= _GEN_4300;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h30 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_48 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h30 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_48 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_48 <= _GEN_4301;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h31 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_49 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h31 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_49 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_49 <= _GEN_4302;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h32 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_50 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h32 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_50 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_50 <= _GEN_4303;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h33 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_51 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h33 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_51 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_51 <= _GEN_4304;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h34 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_52 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h34 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_52 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_52 <= _GEN_4305;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h35 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_53 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h35 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_53 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_53 <= _GEN_4306;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h36 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_54 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h36 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_54 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_54 <= _GEN_4307;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h37 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_55 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h37 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_55 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_55 <= _GEN_4308;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h38 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_56 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h38 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_56 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_56 <= _GEN_4309;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h39 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_57 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h39 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_57 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_57 <= _GEN_4310;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_58 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_58 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_58 <= _GEN_4311;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_59 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_59 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_59 <= _GEN_4312;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_60 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_60 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_60 <= _GEN_4313;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_61 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_61 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_61 <= _GEN_4314;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_62 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_62 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_62 <= _GEN_4315;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_63 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_63 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_63 <= _GEN_4316;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h40 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_64 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h40 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_64 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_64 <= _GEN_4317;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h41 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_65 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h41 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_65 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_65 <= _GEN_4318;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h42 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_66 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h42 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_66 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_66 <= _GEN_4319;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h43 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_67 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h43 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_67 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_67 <= _GEN_4320;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h44 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_68 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h44 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_68 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_68 <= _GEN_4321;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h45 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_69 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h45 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_69 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_69 <= _GEN_4322;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h46 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_70 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h46 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_70 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_70 <= _GEN_4323;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h47 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_71 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h47 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_71 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_71 <= _GEN_4324;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h48 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_72 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h48 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_72 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_72 <= _GEN_4325;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h49 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_73 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h49 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_73 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_73 <= _GEN_4326;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h4a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_74 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h4a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_74 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_74 <= _GEN_4327;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h4b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_75 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h4b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_75 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_75 <= _GEN_4328;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h4c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_76 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h4c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_76 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_76 <= _GEN_4329;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h4d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_77 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h4d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_77 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_77 <= _GEN_4330;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h4e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_78 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h4e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_78 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_78 <= _GEN_4331;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h4f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_79 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h4f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_79 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_79 <= _GEN_4332;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h50 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_80 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h50 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_80 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_80 <= _GEN_4333;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h51 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_81 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h51 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_81 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_81 <= _GEN_4334;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h52 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_82 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h52 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_82 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_82 <= _GEN_4335;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h53 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_83 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h53 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_83 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_83 <= _GEN_4336;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h54 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_84 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h54 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_84 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_84 <= _GEN_4337;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h55 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_85 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h55 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_85 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_85 <= _GEN_4338;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h56 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_86 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h56 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_86 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_86 <= _GEN_4339;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h57 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_87 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h57 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_87 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_87 <= _GEN_4340;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h58 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_88 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h58 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_88 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_88 <= _GEN_4341;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h59 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_89 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h59 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_89 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_89 <= _GEN_4342;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h5a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_90 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h5a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_90 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_90 <= _GEN_4343;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h5b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_91 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h5b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_91 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_91 <= _GEN_4344;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h5c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_92 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h5c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_92 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_92 <= _GEN_4345;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h5d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_93 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h5d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_93 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_93 <= _GEN_4346;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h5e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_94 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h5e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_94 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_94 <= _GEN_4347;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h5f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_95 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h5f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_95 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_95 <= _GEN_4348;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h60 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_96 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h60 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_96 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_96 <= _GEN_4349;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h61 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_97 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h61 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_97 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_97 <= _GEN_4350;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h62 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_98 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h62 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_98 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_98 <= _GEN_4351;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h63 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_99 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h63 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_99 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_99 <= _GEN_4352;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h64 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_100 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h64 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_100 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_100 <= _GEN_4353;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h65 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_101 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h65 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_101 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_101 <= _GEN_4354;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h66 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_102 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h66 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_102 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_102 <= _GEN_4355;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h67 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_103 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h67 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_103 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_103 <= _GEN_4356;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h68 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_104 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h68 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_104 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_104 <= _GEN_4357;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h69 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_105 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h69 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_105 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_105 <= _GEN_4358;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h6a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_106 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h6a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_106 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_106 <= _GEN_4359;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h6b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_107 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h6b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_107 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_107 <= _GEN_4360;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h6c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_108 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h6c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_108 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_108 <= _GEN_4361;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h6d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_109 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h6d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_109 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_109 <= _GEN_4362;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h6e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_110 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h6e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_110 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_110 <= _GEN_4363;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h6f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_111 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h6f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_111 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_111 <= _GEN_4364;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h70 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_112 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h70 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_112 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_112 <= _GEN_4365;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h71 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_113 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h71 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_113 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_113 <= _GEN_4366;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h72 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_114 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h72 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_114 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_114 <= _GEN_4367;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h73 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_115 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h73 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_115 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_115 <= _GEN_4368;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h74 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_116 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h74 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_116 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_116 <= _GEN_4369;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h75 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_117 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h75 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_117 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_117 <= _GEN_4370;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h76 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_118 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h76 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_118 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_118 <= _GEN_4371;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h77 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_119 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h77 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_119 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_119 <= _GEN_4372;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h78 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_120 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h78 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_120 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_120 <= _GEN_4373;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h79 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_121 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h79 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_121 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_121 <= _GEN_4374;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h7a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_122 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h7a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_122 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_122 <= _GEN_4375;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h7b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_123 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h7b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_123 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_123 <= _GEN_4376;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h7c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_124 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h7c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_124 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_124 <= _GEN_4377;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h7d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_125 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h7d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_125 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_125 <= _GEN_4378;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h7e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_126 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h7e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_126 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_126 <= _GEN_4379;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h7f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_127 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h7f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_127 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_127 <= _GEN_4380;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h80 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_128 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h80 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_128 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_128 <= _GEN_4381;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h81 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_129 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h81 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_129 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_129 <= _GEN_4382;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h82 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_130 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h82 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_130 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_130 <= _GEN_4383;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h83 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_131 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h83 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_131 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_131 <= _GEN_4384;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h84 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_132 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h84 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_132 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_132 <= _GEN_4385;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h85 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_133 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h85 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_133 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_133 <= _GEN_4386;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h86 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_134 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h86 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_134 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_134 <= _GEN_4387;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h87 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_135 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h87 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_135 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_135 <= _GEN_4388;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h88 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_136 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h88 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_136 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_136 <= _GEN_4389;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h89 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_137 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h89 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_137 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_137 <= _GEN_4390;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h8a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_138 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h8a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_138 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_138 <= _GEN_4391;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h8b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_139 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h8b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_139 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_139 <= _GEN_4392;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h8c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_140 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h8c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_140 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_140 <= _GEN_4393;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h8d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_141 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h8d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_141 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_141 <= _GEN_4394;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h8e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_142 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h8e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_142 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_142 <= _GEN_4395;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h8f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_143 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h8f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_143 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_143 <= _GEN_4396;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h90 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_144 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h90 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_144 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_144 <= _GEN_4397;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h91 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_145 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h91 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_145 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_145 <= _GEN_4398;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h92 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_146 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h92 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_146 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_146 <= _GEN_4399;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h93 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_147 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h93 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_147 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_147 <= _GEN_4400;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h94 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_148 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h94 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_148 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_148 <= _GEN_4401;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h95 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_149 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h95 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_149 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_149 <= _GEN_4402;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h96 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_150 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h96 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_150 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_150 <= _GEN_4403;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h97 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_151 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h97 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_151 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_151 <= _GEN_4404;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h98 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_152 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h98 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_152 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_152 <= _GEN_4405;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h99 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_153 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h99 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_153 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_153 <= _GEN_4406;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h9a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_154 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h9a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_154 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_154 <= _GEN_4407;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h9b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_155 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h9b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_155 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_155 <= _GEN_4408;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h9c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_156 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h9c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_156 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_156 <= _GEN_4409;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h9d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_157 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h9d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_157 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_157 <= _GEN_4410;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h9e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_158 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h9e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_158 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_158 <= _GEN_4411;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h9f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_159 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h9f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_159 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_159 <= _GEN_4412;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'ha0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_160 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'ha0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_160 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_160 <= _GEN_4413;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'ha1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_161 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'ha1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_161 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_161 <= _GEN_4414;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'ha2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_162 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'ha2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_162 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_162 <= _GEN_4415;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'ha3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_163 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'ha3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_163 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_163 <= _GEN_4416;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'ha4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_164 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'ha4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_164 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_164 <= _GEN_4417;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'ha5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_165 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'ha5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_165 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_165 <= _GEN_4418;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'ha6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_166 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'ha6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_166 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_166 <= _GEN_4419;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'ha7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_167 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'ha7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_167 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_167 <= _GEN_4420;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'ha8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_168 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'ha8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_168 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_168 <= _GEN_4421;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'ha9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_169 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'ha9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_169 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_169 <= _GEN_4422;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'haa == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_170 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'haa == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_170 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_170 <= _GEN_4423;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hab == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_171 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hab == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_171 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_171 <= _GEN_4424;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hac == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_172 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hac == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_172 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_172 <= _GEN_4425;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'had == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_173 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'had == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_173 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_173 <= _GEN_4426;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hae == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_174 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hae == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_174 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_174 <= _GEN_4427;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'haf == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_175 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'haf == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_175 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_175 <= _GEN_4428;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hb0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_176 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hb0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_176 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_176 <= _GEN_4429;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hb1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_177 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hb1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_177 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_177 <= _GEN_4430;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hb2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_178 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hb2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_178 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_178 <= _GEN_4431;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hb3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_179 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hb3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_179 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_179 <= _GEN_4432;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hb4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_180 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hb4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_180 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_180 <= _GEN_4433;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hb5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_181 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hb5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_181 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_181 <= _GEN_4434;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hb6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_182 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hb6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_182 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_182 <= _GEN_4435;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hb7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_183 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hb7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_183 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_183 <= _GEN_4436;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hb8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_184 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hb8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_184 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_184 <= _GEN_4437;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hb9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_185 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hb9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_185 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_185 <= _GEN_4438;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hba == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_186 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hba == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_186 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_186 <= _GEN_4439;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hbb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_187 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hbb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_187 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_187 <= _GEN_4440;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hbc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_188 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hbc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_188 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_188 <= _GEN_4441;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hbd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_189 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hbd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_189 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_189 <= _GEN_4442;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hbe == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_190 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hbe == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_190 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_190 <= _GEN_4443;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hbf == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_191 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hbf == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_191 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_191 <= _GEN_4444;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hc0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_192 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hc0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_192 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_192 <= _GEN_4445;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hc1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_193 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hc1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_193 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_193 <= _GEN_4446;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hc2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_194 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hc2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_194 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_194 <= _GEN_4447;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hc3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_195 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hc3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_195 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_195 <= _GEN_4448;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hc4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_196 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hc4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_196 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_196 <= _GEN_4449;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hc5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_197 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hc5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_197 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_197 <= _GEN_4450;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hc6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_198 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hc6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_198 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_198 <= _GEN_4451;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hc7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_199 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hc7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_199 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_199 <= _GEN_4452;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hc8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_200 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hc8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_200 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_200 <= _GEN_4453;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hc9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_201 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hc9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_201 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_201 <= _GEN_4454;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hca == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_202 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hca == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_202 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_202 <= _GEN_4455;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hcb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_203 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hcb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_203 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_203 <= _GEN_4456;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hcc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_204 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hcc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_204 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_204 <= _GEN_4457;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hcd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_205 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hcd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_205 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_205 <= _GEN_4458;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hce == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_206 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hce == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_206 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_206 <= _GEN_4459;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hcf == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_207 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hcf == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_207 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_207 <= _GEN_4460;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hd0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_208 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hd0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_208 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_208 <= _GEN_4461;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hd1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_209 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hd1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_209 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_209 <= _GEN_4462;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hd2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_210 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hd2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_210 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_210 <= _GEN_4463;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hd3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_211 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hd3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_211 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_211 <= _GEN_4464;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hd4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_212 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hd4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_212 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_212 <= _GEN_4465;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hd5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_213 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hd5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_213 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_213 <= _GEN_4466;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hd6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_214 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hd6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_214 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_214 <= _GEN_4467;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hd7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_215 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hd7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_215 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_215 <= _GEN_4468;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hd8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_216 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hd8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_216 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_216 <= _GEN_4469;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hd9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_217 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hd9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_217 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_217 <= _GEN_4470;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hda == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_218 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hda == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_218 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_218 <= _GEN_4471;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hdb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_219 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hdb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_219 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_219 <= _GEN_4472;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hdc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_220 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hdc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_220 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_220 <= _GEN_4473;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hdd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_221 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hdd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_221 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_221 <= _GEN_4474;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hde == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_222 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hde == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_222 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_222 <= _GEN_4475;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hdf == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_223 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hdf == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_223 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_223 <= _GEN_4476;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'he0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_224 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'he0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_224 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_224 <= _GEN_4477;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'he1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_225 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'he1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_225 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_225 <= _GEN_4478;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'he2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_226 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'he2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_226 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_226 <= _GEN_4479;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'he3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_227 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'he3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_227 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_227 <= _GEN_4480;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'he4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_228 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'he4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_228 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_228 <= _GEN_4481;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'he5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_229 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'he5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_229 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_229 <= _GEN_4482;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'he6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_230 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'he6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_230 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_230 <= _GEN_4483;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'he7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_231 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'he7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_231 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_231 <= _GEN_4484;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'he8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_232 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'he8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_232 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_232 <= _GEN_4485;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'he9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_233 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'he9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_233 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_233 <= _GEN_4486;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hea == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_234 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hea == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_234 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_234 <= _GEN_4487;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'heb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_235 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'heb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_235 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_235 <= _GEN_4488;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hec == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_236 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hec == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_236 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_236 <= _GEN_4489;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hed == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_237 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hed == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_237 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_237 <= _GEN_4490;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hee == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_238 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hee == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_238 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_238 <= _GEN_4491;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hef == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_239 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hef == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_239 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_239 <= _GEN_4492;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hf0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_240 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hf0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_240 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_240 <= _GEN_4493;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hf1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_241 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hf1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_241 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_241 <= _GEN_4494;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hf2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_242 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hf2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_242 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_242 <= _GEN_4495;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hf3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_243 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hf3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_243 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_243 <= _GEN_4496;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hf4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_244 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hf4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_244 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_244 <= _GEN_4497;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hf5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_245 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hf5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_245 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_245 <= _GEN_4498;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hf6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_246 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hf6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_246 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_246 <= _GEN_4499;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hf7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_247 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hf7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_247 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_247 <= _GEN_4500;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hf8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_248 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hf8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_248 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_248 <= _GEN_4501;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hf9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_249 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hf9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_249 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_249 <= _GEN_4502;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hfa == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_250 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hfa == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_250 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_250 <= _GEN_4503;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hfb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_251 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hfb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_251 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_251 <= _GEN_4504;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hfc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_252 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hfc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_252 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_252 <= _GEN_4505;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hfd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_253 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hfd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_253 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_253 <= _GEN_4506;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hfe == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_254 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hfe == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_254 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_254 <= _GEN_4507;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'hff == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_255 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'hff == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_255 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_255 <= _GEN_4508;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h100 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_256 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h100 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_256 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_256 <= _GEN_4509;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h101 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_257 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h101 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_257 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_257 <= _GEN_4510;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h102 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_258 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h102 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_258 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_258 <= _GEN_4511;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h103 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_259 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h103 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_259 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_259 <= _GEN_4512;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h104 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_260 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h104 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_260 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_260 <= _GEN_4513;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h105 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_261 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h105 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_261 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_261 <= _GEN_4514;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h106 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_262 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h106 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_262 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_262 <= _GEN_4515;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h107 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_263 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h107 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_263 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_263 <= _GEN_4516;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h108 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_264 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h108 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_264 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_264 <= _GEN_4517;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h109 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_265 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h109 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_265 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_265 <= _GEN_4518;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h10a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_266 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h10a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_266 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_266 <= _GEN_4519;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h10b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_267 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h10b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_267 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_267 <= _GEN_4520;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h10c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_268 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h10c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_268 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_268 <= _GEN_4521;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h10d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_269 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h10d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_269 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_269 <= _GEN_4522;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h10e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_270 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h10e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_270 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_270 <= _GEN_4523;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h10f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_271 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h10f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_271 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_271 <= _GEN_4524;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h110 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_272 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h110 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_272 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_272 <= _GEN_4525;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h111 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_273 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h111 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_273 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_273 <= _GEN_4526;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h112 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_274 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h112 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_274 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_274 <= _GEN_4527;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h113 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_275 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h113 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_275 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_275 <= _GEN_4528;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h114 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_276 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h114 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_276 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_276 <= _GEN_4529;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h115 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_277 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h115 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_277 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_277 <= _GEN_4530;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h116 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_278 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h116 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_278 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_278 <= _GEN_4531;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h117 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_279 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h117 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_279 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_279 <= _GEN_4532;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h118 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_280 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h118 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_280 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_280 <= _GEN_4533;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h119 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_281 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h119 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_281 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_281 <= _GEN_4534;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h11a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_282 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h11a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_282 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_282 <= _GEN_4535;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h11b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_283 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h11b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_283 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_283 <= _GEN_4536;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h11c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_284 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h11c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_284 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_284 <= _GEN_4537;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h11d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_285 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h11d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_285 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_285 <= _GEN_4538;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h11e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_286 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h11e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_286 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_286 <= _GEN_4539;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h11f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_287 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h11f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_287 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_287 <= _GEN_4540;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h120 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_288 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h120 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_288 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_288 <= _GEN_4541;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h121 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_289 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h121 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_289 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_289 <= _GEN_4542;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h122 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_290 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h122 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_290 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_290 <= _GEN_4543;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h123 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_291 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h123 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_291 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_291 <= _GEN_4544;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h124 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_292 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h124 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_292 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_292 <= _GEN_4545;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h125 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_293 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h125 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_293 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_293 <= _GEN_4546;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h126 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_294 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h126 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_294 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_294 <= _GEN_4547;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h127 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_295 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h127 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_295 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_295 <= _GEN_4548;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h128 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_296 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h128 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_296 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_296 <= _GEN_4549;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h129 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_297 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h129 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_297 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_297 <= _GEN_4550;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h12a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_298 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h12a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_298 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_298 <= _GEN_4551;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h12b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_299 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h12b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_299 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_299 <= _GEN_4552;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h12c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_300 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h12c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_300 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_300 <= _GEN_4553;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h12d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_301 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h12d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_301 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_301 <= _GEN_4554;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h12e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_302 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h12e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_302 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_302 <= _GEN_4555;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h12f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_303 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h12f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_303 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_303 <= _GEN_4556;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h130 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_304 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h130 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_304 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_304 <= _GEN_4557;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h131 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_305 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h131 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_305 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_305 <= _GEN_4558;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h132 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_306 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h132 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_306 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_306 <= _GEN_4559;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h133 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_307 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h133 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_307 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_307 <= _GEN_4560;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h134 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_308 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h134 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_308 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_308 <= _GEN_4561;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h135 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_309 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h135 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_309 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_309 <= _GEN_4562;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h136 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_310 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h136 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_310 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_310 <= _GEN_4563;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h137 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_311 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h137 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_311 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_311 <= _GEN_4564;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h138 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_312 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h138 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_312 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_312 <= _GEN_4565;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h139 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_313 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h139 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_313 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_313 <= _GEN_4566;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h13a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_314 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h13a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_314 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_314 <= _GEN_4567;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h13b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_315 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h13b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_315 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_315 <= _GEN_4568;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h13c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_316 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h13c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_316 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_316 <= _GEN_4569;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h13d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_317 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h13d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_317 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_317 <= _GEN_4570;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h13e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_318 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h13e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_318 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_318 <= _GEN_4571;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h13f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_319 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h13f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_319 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_319 <= _GEN_4572;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h140 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_320 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h140 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_320 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_320 <= _GEN_4573;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h141 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_321 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h141 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_321 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_321 <= _GEN_4574;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h142 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_322 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h142 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_322 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_322 <= _GEN_4575;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h143 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_323 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h143 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_323 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_323 <= _GEN_4576;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h144 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_324 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h144 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_324 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_324 <= _GEN_4577;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h145 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_325 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h145 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_325 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_325 <= _GEN_4578;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h146 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_326 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h146 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_326 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_326 <= _GEN_4579;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h147 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_327 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h147 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_327 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_327 <= _GEN_4580;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h148 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_328 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h148 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_328 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_328 <= _GEN_4581;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h149 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_329 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h149 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_329 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_329 <= _GEN_4582;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h14a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_330 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h14a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_330 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_330 <= _GEN_4583;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h14b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_331 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h14b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_331 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_331 <= _GEN_4584;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h14c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_332 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h14c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_332 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_332 <= _GEN_4585;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h14d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_333 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h14d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_333 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_333 <= _GEN_4586;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h14e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_334 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h14e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_334 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_334 <= _GEN_4587;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h14f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_335 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h14f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_335 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_335 <= _GEN_4588;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h150 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_336 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h150 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_336 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_336 <= _GEN_4589;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h151 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_337 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h151 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_337 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_337 <= _GEN_4590;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h152 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_338 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h152 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_338 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_338 <= _GEN_4591;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h153 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_339 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h153 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_339 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_339 <= _GEN_4592;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h154 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_340 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h154 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_340 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_340 <= _GEN_4593;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h155 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_341 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h155 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_341 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_341 <= _GEN_4594;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h156 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_342 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h156 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_342 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_342 <= _GEN_4595;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h157 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_343 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h157 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_343 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_343 <= _GEN_4596;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h158 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_344 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h158 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_344 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_344 <= _GEN_4597;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h159 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_345 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h159 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_345 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_345 <= _GEN_4598;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h15a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_346 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h15a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_346 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_346 <= _GEN_4599;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h15b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_347 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h15b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_347 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_347 <= _GEN_4600;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h15c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_348 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h15c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_348 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_348 <= _GEN_4601;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h15d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_349 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h15d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_349 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_349 <= _GEN_4602;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h15e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_350 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h15e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_350 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_350 <= _GEN_4603;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h15f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_351 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h15f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_351 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_351 <= _GEN_4604;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h160 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_352 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h160 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_352 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_352 <= _GEN_4605;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h161 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_353 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h161 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_353 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_353 <= _GEN_4606;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h162 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_354 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h162 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_354 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_354 <= _GEN_4607;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h163 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_355 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h163 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_355 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_355 <= _GEN_4608;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h164 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_356 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h164 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_356 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_356 <= _GEN_4609;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h165 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_357 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h165 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_357 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_357 <= _GEN_4610;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h166 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_358 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h166 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_358 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_358 <= _GEN_4611;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h167 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_359 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h167 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_359 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_359 <= _GEN_4612;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h168 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_360 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h168 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_360 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_360 <= _GEN_4613;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h169 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_361 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h169 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_361 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_361 <= _GEN_4614;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h16a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_362 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h16a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_362 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_362 <= _GEN_4615;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h16b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_363 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h16b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_363 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_363 <= _GEN_4616;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h16c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_364 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h16c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_364 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_364 <= _GEN_4617;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h16d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_365 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h16d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_365 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_365 <= _GEN_4618;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h16e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_366 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h16e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_366 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_366 <= _GEN_4619;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h16f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_367 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h16f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_367 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_367 <= _GEN_4620;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h170 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_368 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h170 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_368 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_368 <= _GEN_4621;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h171 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_369 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h171 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_369 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_369 <= _GEN_4622;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h172 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_370 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h172 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_370 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_370 <= _GEN_4623;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h173 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_371 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h173 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_371 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_371 <= _GEN_4624;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h174 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_372 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h174 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_372 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_372 <= _GEN_4625;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h175 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_373 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h175 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_373 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_373 <= _GEN_4626;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h176 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_374 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h176 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_374 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_374 <= _GEN_4627;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h177 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_375 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h177 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_375 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_375 <= _GEN_4628;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h178 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_376 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h178 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_376 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_376 <= _GEN_4629;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h179 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_377 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h179 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_377 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_377 <= _GEN_4630;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h17a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_378 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h17a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_378 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_378 <= _GEN_4631;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h17b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_379 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h17b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_379 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_379 <= _GEN_4632;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h17c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_380 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h17c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_380 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_380 <= _GEN_4633;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h17d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_381 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h17d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_381 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_381 <= _GEN_4634;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h17e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_382 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h17e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_382 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_382 <= _GEN_4635;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h17f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_383 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h17f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_383 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_383 <= _GEN_4636;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h180 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_384 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h180 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_384 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_384 <= _GEN_4637;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h181 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_385 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h181 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_385 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_385 <= _GEN_4638;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h182 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_386 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h182 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_386 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_386 <= _GEN_4639;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h183 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_387 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h183 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_387 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_387 <= _GEN_4640;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h184 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_388 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h184 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_388 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_388 <= _GEN_4641;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h185 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_389 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h185 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_389 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_389 <= _GEN_4642;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h186 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_390 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h186 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_390 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_390 <= _GEN_4643;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h187 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_391 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h187 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_391 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_391 <= _GEN_4644;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h188 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_392 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h188 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_392 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_392 <= _GEN_4645;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h189 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_393 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h189 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_393 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_393 <= _GEN_4646;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h18a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_394 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h18a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_394 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_394 <= _GEN_4647;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h18b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_395 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h18b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_395 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_395 <= _GEN_4648;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h18c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_396 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h18c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_396 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_396 <= _GEN_4649;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h18d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_397 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h18d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_397 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_397 <= _GEN_4650;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h18e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_398 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h18e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_398 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_398 <= _GEN_4651;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h18f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_399 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h18f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_399 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_399 <= _GEN_4652;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h190 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_400 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h190 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_400 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_400 <= _GEN_4653;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h191 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_401 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h191 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_401 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_401 <= _GEN_4654;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h192 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_402 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h192 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_402 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_402 <= _GEN_4655;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h193 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_403 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h193 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_403 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_403 <= _GEN_4656;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h194 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_404 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h194 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_404 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_404 <= _GEN_4657;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h195 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_405 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h195 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_405 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_405 <= _GEN_4658;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h196 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_406 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h196 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_406 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_406 <= _GEN_4659;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h197 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_407 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h197 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_407 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_407 <= _GEN_4660;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h198 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_408 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h198 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_408 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_408 <= _GEN_4661;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h199 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_409 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h199 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_409 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_409 <= _GEN_4662;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h19a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_410 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h19a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_410 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_410 <= _GEN_4663;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h19b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_411 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h19b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_411 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_411 <= _GEN_4664;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h19c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_412 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h19c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_412 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_412 <= _GEN_4665;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h19d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_413 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h19d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_413 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_413 <= _GEN_4666;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h19e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_414 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h19e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_414 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_414 <= _GEN_4667;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h19f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_415 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h19f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_415 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_415 <= _GEN_4668;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1a0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_416 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1a0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_416 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_416 <= _GEN_4669;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1a1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_417 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1a1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_417 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_417 <= _GEN_4670;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1a2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_418 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1a2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_418 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_418 <= _GEN_4671;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1a3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_419 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1a3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_419 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_419 <= _GEN_4672;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1a4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_420 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1a4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_420 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_420 <= _GEN_4673;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1a5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_421 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1a5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_421 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_421 <= _GEN_4674;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1a6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_422 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1a6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_422 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_422 <= _GEN_4675;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1a7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_423 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1a7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_423 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_423 <= _GEN_4676;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1a8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_424 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1a8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_424 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_424 <= _GEN_4677;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1a9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_425 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1a9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_425 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_425 <= _GEN_4678;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1aa == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_426 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1aa == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_426 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_426 <= _GEN_4679;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ab == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_427 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ab == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_427 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_427 <= _GEN_4680;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ac == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_428 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ac == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_428 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_428 <= _GEN_4681;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ad == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_429 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ad == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_429 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_429 <= _GEN_4682;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ae == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_430 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ae == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_430 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_430 <= _GEN_4683;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1af == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_431 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1af == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_431 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_431 <= _GEN_4684;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1b0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_432 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1b0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_432 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_432 <= _GEN_4685;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1b1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_433 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1b1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_433 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_433 <= _GEN_4686;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1b2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_434 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1b2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_434 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_434 <= _GEN_4687;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1b3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_435 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1b3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_435 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_435 <= _GEN_4688;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1b4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_436 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1b4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_436 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_436 <= _GEN_4689;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1b5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_437 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1b5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_437 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_437 <= _GEN_4690;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1b6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_438 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1b6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_438 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_438 <= _GEN_4691;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1b7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_439 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1b7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_439 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_439 <= _GEN_4692;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1b8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_440 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1b8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_440 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_440 <= _GEN_4693;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1b9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_441 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1b9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_441 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_441 <= _GEN_4694;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ba == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_442 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ba == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_442 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_442 <= _GEN_4695;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1bb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_443 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1bb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_443 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_443 <= _GEN_4696;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1bc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_444 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1bc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_444 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_444 <= _GEN_4697;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1bd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_445 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1bd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_445 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_445 <= _GEN_4698;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1be == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_446 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1be == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_446 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_446 <= _GEN_4699;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1bf == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_447 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1bf == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_447 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_447 <= _GEN_4700;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1c0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_448 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1c0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_448 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_448 <= _GEN_4701;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1c1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_449 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1c1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_449 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_449 <= _GEN_4702;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1c2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_450 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1c2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_450 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_450 <= _GEN_4703;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1c3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_451 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1c3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_451 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_451 <= _GEN_4704;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1c4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_452 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1c4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_452 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_452 <= _GEN_4705;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1c5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_453 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1c5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_453 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_453 <= _GEN_4706;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1c6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_454 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1c6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_454 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_454 <= _GEN_4707;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1c7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_455 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1c7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_455 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_455 <= _GEN_4708;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1c8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_456 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1c8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_456 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_456 <= _GEN_4709;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1c9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_457 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1c9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_457 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_457 <= _GEN_4710;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ca == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_458 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ca == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_458 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_458 <= _GEN_4711;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1cb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_459 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1cb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_459 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_459 <= _GEN_4712;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1cc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_460 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1cc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_460 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_460 <= _GEN_4713;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1cd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_461 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1cd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_461 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_461 <= _GEN_4714;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ce == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_462 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ce == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_462 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_462 <= _GEN_4715;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1cf == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_463 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1cf == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_463 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_463 <= _GEN_4716;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1d0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_464 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1d0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_464 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_464 <= _GEN_4717;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1d1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_465 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1d1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_465 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_465 <= _GEN_4718;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1d2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_466 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1d2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_466 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_466 <= _GEN_4719;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1d3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_467 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1d3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_467 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_467 <= _GEN_4720;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1d4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_468 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1d4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_468 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_468 <= _GEN_4721;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1d5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_469 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1d5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_469 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_469 <= _GEN_4722;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1d6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_470 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1d6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_470 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_470 <= _GEN_4723;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1d7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_471 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1d7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_471 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_471 <= _GEN_4724;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1d8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_472 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1d8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_472 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_472 <= _GEN_4725;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1d9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_473 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1d9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_473 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_473 <= _GEN_4726;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1da == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_474 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1da == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_474 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_474 <= _GEN_4727;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1db == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_475 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1db == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_475 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_475 <= _GEN_4728;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1dc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_476 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1dc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_476 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_476 <= _GEN_4729;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1dd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_477 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1dd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_477 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_477 <= _GEN_4730;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1de == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_478 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1de == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_478 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_478 <= _GEN_4731;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1df == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_479 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1df == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_479 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_479 <= _GEN_4732;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1e0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_480 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1e0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_480 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_480 <= _GEN_4733;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1e1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_481 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1e1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_481 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_481 <= _GEN_4734;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1e2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_482 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1e2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_482 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_482 <= _GEN_4735;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1e3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_483 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1e3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_483 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_483 <= _GEN_4736;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1e4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_484 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1e4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_484 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_484 <= _GEN_4737;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1e5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_485 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1e5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_485 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_485 <= _GEN_4738;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1e6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_486 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1e6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_486 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_486 <= _GEN_4739;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1e7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_487 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1e7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_487 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_487 <= _GEN_4740;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1e8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_488 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1e8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_488 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_488 <= _GEN_4741;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1e9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_489 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1e9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_489 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_489 <= _GEN_4742;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ea == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_490 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ea == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_490 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_490 <= _GEN_4743;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1eb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_491 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1eb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_491 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_491 <= _GEN_4744;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ec == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_492 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ec == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_492 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_492 <= _GEN_4745;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ed == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_493 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ed == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_493 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_493 <= _GEN_4746;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ee == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_494 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ee == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_494 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_494 <= _GEN_4747;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ef == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_495 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ef == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_495 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_495 <= _GEN_4748;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1f0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_496 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1f0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_496 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_496 <= _GEN_4749;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1f1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_497 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1f1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_497 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_497 <= _GEN_4750;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1f2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_498 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1f2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_498 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_498 <= _GEN_4751;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1f3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_499 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1f3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_499 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_499 <= _GEN_4752;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1f4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_500 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1f4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_500 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_500 <= _GEN_4753;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1f5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_501 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1f5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_501 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_501 <= _GEN_4754;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1f6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_502 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1f6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_502 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_502 <= _GEN_4755;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1f7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_503 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1f7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_503 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_503 <= _GEN_4756;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1f8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_504 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1f8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_504 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_504 <= _GEN_4757;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1f9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_505 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1f9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_505 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_505 <= _GEN_4758;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1fa == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_506 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1fa == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_506 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_506 <= _GEN_4759;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1fb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_507 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1fb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_507 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_507 <= _GEN_4760;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1fc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_508 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1fc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_508 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_508 <= _GEN_4761;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1fd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_509 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1fd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_509 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_509 <= _GEN_4762;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1fe == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_510 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1fe == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_510 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_510 <= _GEN_4763;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h1ff == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_511 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h1ff == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_511 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_511 <= _GEN_4764;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h200 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_512 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h200 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_512 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_512 <= _GEN_4765;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h201 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_513 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h201 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_513 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_513 <= _GEN_4766;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h202 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_514 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h202 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_514 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_514 <= _GEN_4767;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h203 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_515 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h203 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_515 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_515 <= _GEN_4768;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h204 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_516 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h204 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_516 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_516 <= _GEN_4769;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h205 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_517 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h205 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_517 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_517 <= _GEN_4770;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h206 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_518 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h206 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_518 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_518 <= _GEN_4771;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h207 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_519 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h207 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_519 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_519 <= _GEN_4772;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h208 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_520 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h208 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_520 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_520 <= _GEN_4773;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h209 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_521 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h209 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_521 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_521 <= _GEN_4774;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h20a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_522 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h20a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_522 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_522 <= _GEN_4775;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h20b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_523 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h20b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_523 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_523 <= _GEN_4776;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h20c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_524 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h20c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_524 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_524 <= _GEN_4777;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h20d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_525 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h20d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_525 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_525 <= _GEN_4778;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h20e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_526 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h20e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_526 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_526 <= _GEN_4779;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h20f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_527 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h20f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_527 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_527 <= _GEN_4780;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h210 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_528 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h210 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_528 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_528 <= _GEN_4781;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h211 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_529 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h211 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_529 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_529 <= _GEN_4782;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h212 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_530 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h212 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_530 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_530 <= _GEN_4783;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h213 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_531 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h213 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_531 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_531 <= _GEN_4784;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h214 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_532 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h214 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_532 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_532 <= _GEN_4785;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h215 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_533 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h215 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_533 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_533 <= _GEN_4786;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h216 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_534 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h216 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_534 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_534 <= _GEN_4787;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h217 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_535 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h217 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_535 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_535 <= _GEN_4788;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h218 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_536 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h218 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_536 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_536 <= _GEN_4789;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h219 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_537 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h219 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_537 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_537 <= _GEN_4790;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h21a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_538 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h21a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_538 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_538 <= _GEN_4791;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h21b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_539 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h21b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_539 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_539 <= _GEN_4792;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h21c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_540 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h21c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_540 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_540 <= _GEN_4793;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h21d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_541 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h21d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_541 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_541 <= _GEN_4794;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h21e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_542 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h21e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_542 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_542 <= _GEN_4795;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h21f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_543 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h21f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_543 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_543 <= _GEN_4796;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h220 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_544 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h220 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_544 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_544 <= _GEN_4797;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h221 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_545 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h221 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_545 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_545 <= _GEN_4798;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h222 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_546 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h222 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_546 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_546 <= _GEN_4799;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h223 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_547 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h223 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_547 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_547 <= _GEN_4800;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h224 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_548 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h224 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_548 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_548 <= _GEN_4801;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h225 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_549 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h225 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_549 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_549 <= _GEN_4802;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h226 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_550 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h226 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_550 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_550 <= _GEN_4803;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h227 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_551 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h227 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_551 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_551 <= _GEN_4804;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h228 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_552 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h228 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_552 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_552 <= _GEN_4805;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h229 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_553 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h229 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_553 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_553 <= _GEN_4806;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h22a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_554 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h22a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_554 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_554 <= _GEN_4807;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h22b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_555 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h22b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_555 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_555 <= _GEN_4808;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h22c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_556 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h22c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_556 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_556 <= _GEN_4809;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h22d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_557 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h22d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_557 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_557 <= _GEN_4810;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h22e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_558 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h22e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_558 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_558 <= _GEN_4811;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h22f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_559 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h22f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_559 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_559 <= _GEN_4812;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h230 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_560 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h230 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_560 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_560 <= _GEN_4813;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h231 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_561 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h231 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_561 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_561 <= _GEN_4814;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h232 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_562 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h232 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_562 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_562 <= _GEN_4815;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h233 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_563 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h233 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_563 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_563 <= _GEN_4816;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h234 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_564 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h234 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_564 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_564 <= _GEN_4817;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h235 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_565 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h235 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_565 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_565 <= _GEN_4818;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h236 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_566 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h236 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_566 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_566 <= _GEN_4819;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h237 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_567 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h237 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_567 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_567 <= _GEN_4820;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h238 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_568 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h238 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_568 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_568 <= _GEN_4821;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h239 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_569 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h239 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_569 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_569 <= _GEN_4822;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h23a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_570 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h23a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_570 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_570 <= _GEN_4823;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h23b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_571 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h23b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_571 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_571 <= _GEN_4824;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h23c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_572 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h23c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_572 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_572 <= _GEN_4825;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h23d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_573 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h23d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_573 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_573 <= _GEN_4826;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h23e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_574 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h23e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_574 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_574 <= _GEN_4827;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h23f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_575 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h23f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_575 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_575 <= _GEN_4828;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h240 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_576 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h240 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_576 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_576 <= _GEN_4829;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h241 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_577 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h241 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_577 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_577 <= _GEN_4830;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h242 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_578 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h242 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_578 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_578 <= _GEN_4831;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h243 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_579 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h243 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_579 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_579 <= _GEN_4832;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h244 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_580 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h244 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_580 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_580 <= _GEN_4833;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h245 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_581 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h245 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_581 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_581 <= _GEN_4834;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h246 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_582 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h246 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_582 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_582 <= _GEN_4835;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h247 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_583 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h247 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_583 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_583 <= _GEN_4836;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h248 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_584 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h248 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_584 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_584 <= _GEN_4837;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h249 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_585 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h249 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_585 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_585 <= _GEN_4838;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h24a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_586 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h24a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_586 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_586 <= _GEN_4839;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h24b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_587 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h24b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_587 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_587 <= _GEN_4840;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h24c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_588 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h24c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_588 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_588 <= _GEN_4841;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h24d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_589 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h24d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_589 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_589 <= _GEN_4842;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h24e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_590 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h24e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_590 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_590 <= _GEN_4843;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h24f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_591 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h24f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_591 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_591 <= _GEN_4844;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h250 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_592 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h250 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_592 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_592 <= _GEN_4845;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h251 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_593 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h251 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_593 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_593 <= _GEN_4846;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h252 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_594 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h252 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_594 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_594 <= _GEN_4847;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h253 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_595 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h253 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_595 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_595 <= _GEN_4848;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h254 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_596 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h254 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_596 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_596 <= _GEN_4849;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h255 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_597 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h255 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_597 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_597 <= _GEN_4850;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h256 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_598 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h256 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_598 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_598 <= _GEN_4851;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h257 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_599 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h257 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_599 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_599 <= _GEN_4852;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h258 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_600 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h258 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_600 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_600 <= _GEN_4853;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h259 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_601 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h259 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_601 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_601 <= _GEN_4854;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h25a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_602 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h25a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_602 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_602 <= _GEN_4855;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h25b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_603 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h25b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_603 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_603 <= _GEN_4856;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h25c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_604 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h25c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_604 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_604 <= _GEN_4857;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h25d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_605 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h25d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_605 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_605 <= _GEN_4858;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h25e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_606 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h25e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_606 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_606 <= _GEN_4859;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h25f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_607 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h25f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_607 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_607 <= _GEN_4860;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h260 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_608 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h260 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_608 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_608 <= _GEN_4861;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h261 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_609 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h261 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_609 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_609 <= _GEN_4862;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h262 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_610 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h262 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_610 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_610 <= _GEN_4863;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h263 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_611 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h263 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_611 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_611 <= _GEN_4864;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h264 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_612 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h264 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_612 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_612 <= _GEN_4865;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h265 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_613 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h265 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_613 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_613 <= _GEN_4866;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h266 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_614 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h266 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_614 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_614 <= _GEN_4867;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h267 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_615 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h267 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_615 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_615 <= _GEN_4868;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h268 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_616 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h268 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_616 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_616 <= _GEN_4869;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h269 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_617 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h269 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_617 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_617 <= _GEN_4870;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h26a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_618 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h26a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_618 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_618 <= _GEN_4871;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h26b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_619 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h26b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_619 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_619 <= _GEN_4872;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h26c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_620 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h26c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_620 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_620 <= _GEN_4873;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h26d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_621 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h26d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_621 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_621 <= _GEN_4874;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h26e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_622 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h26e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_622 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_622 <= _GEN_4875;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h26f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_623 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h26f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_623 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_623 <= _GEN_4876;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h270 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_624 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h270 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_624 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_624 <= _GEN_4877;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h271 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_625 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h271 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_625 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_625 <= _GEN_4878;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h272 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_626 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h272 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_626 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_626 <= _GEN_4879;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h273 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_627 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h273 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_627 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_627 <= _GEN_4880;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h274 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_628 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h274 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_628 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_628 <= _GEN_4881;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h275 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_629 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h275 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_629 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_629 <= _GEN_4882;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h276 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_630 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h276 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_630 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_630 <= _GEN_4883;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h277 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_631 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h277 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_631 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_631 <= _GEN_4884;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h278 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_632 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h278 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_632 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_632 <= _GEN_4885;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h279 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_633 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h279 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_633 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_633 <= _GEN_4886;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h27a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_634 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h27a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_634 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_634 <= _GEN_4887;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h27b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_635 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h27b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_635 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_635 <= _GEN_4888;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h27c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_636 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h27c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_636 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_636 <= _GEN_4889;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h27d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_637 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h27d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_637 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_637 <= _GEN_4890;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h27e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_638 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h27e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_638 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_638 <= _GEN_4891;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h27f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_639 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h27f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_639 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_639 <= _GEN_4892;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h280 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_640 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h280 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_640 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_640 <= _GEN_4893;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h281 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_641 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h281 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_641 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_641 <= _GEN_4894;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h282 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_642 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h282 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_642 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_642 <= _GEN_4895;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h283 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_643 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h283 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_643 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_643 <= _GEN_4896;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h284 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_644 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h284 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_644 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_644 <= _GEN_4897;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h285 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_645 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h285 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_645 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_645 <= _GEN_4898;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h286 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_646 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h286 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_646 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_646 <= _GEN_4899;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h287 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_647 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h287 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_647 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_647 <= _GEN_4900;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h288 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_648 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h288 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_648 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_648 <= _GEN_4901;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h289 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_649 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h289 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_649 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_649 <= _GEN_4902;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h28a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_650 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h28a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_650 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_650 <= _GEN_4903;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h28b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_651 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h28b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_651 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_651 <= _GEN_4904;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h28c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_652 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h28c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_652 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_652 <= _GEN_4905;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h28d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_653 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h28d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_653 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_653 <= _GEN_4906;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h28e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_654 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h28e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_654 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_654 <= _GEN_4907;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h28f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_655 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h28f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_655 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_655 <= _GEN_4908;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h290 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_656 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h290 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_656 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_656 <= _GEN_4909;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h291 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_657 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h291 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_657 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_657 <= _GEN_4910;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h292 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_658 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h292 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_658 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_658 <= _GEN_4911;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h293 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_659 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h293 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_659 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_659 <= _GEN_4912;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h294 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_660 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h294 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_660 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_660 <= _GEN_4913;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h295 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_661 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h295 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_661 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_661 <= _GEN_4914;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h296 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_662 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h296 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_662 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_662 <= _GEN_4915;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h297 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_663 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h297 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_663 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_663 <= _GEN_4916;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h298 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_664 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h298 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_664 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_664 <= _GEN_4917;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h299 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_665 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h299 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_665 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_665 <= _GEN_4918;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h29a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_666 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h29a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_666 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_666 <= _GEN_4919;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h29b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_667 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h29b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_667 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_667 <= _GEN_4920;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h29c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_668 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h29c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_668 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_668 <= _GEN_4921;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h29d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_669 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h29d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_669 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_669 <= _GEN_4922;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h29e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_670 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h29e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_670 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_670 <= _GEN_4923;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h29f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_671 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h29f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_671 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_671 <= _GEN_4924;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2a0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_672 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2a0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_672 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_672 <= _GEN_4925;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2a1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_673 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2a1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_673 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_673 <= _GEN_4926;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2a2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_674 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2a2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_674 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_674 <= _GEN_4927;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2a3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_675 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2a3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_675 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_675 <= _GEN_4928;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2a4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_676 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2a4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_676 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_676 <= _GEN_4929;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2a5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_677 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2a5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_677 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_677 <= _GEN_4930;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2a6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_678 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2a6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_678 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_678 <= _GEN_4931;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2a7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_679 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2a7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_679 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_679 <= _GEN_4932;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2a8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_680 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2a8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_680 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_680 <= _GEN_4933;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2a9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_681 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2a9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_681 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_681 <= _GEN_4934;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2aa == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_682 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2aa == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_682 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_682 <= _GEN_4935;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ab == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_683 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ab == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_683 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_683 <= _GEN_4936;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ac == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_684 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ac == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_684 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_684 <= _GEN_4937;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ad == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_685 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ad == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_685 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_685 <= _GEN_4938;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ae == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_686 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ae == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_686 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_686 <= _GEN_4939;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2af == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_687 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2af == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_687 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_687 <= _GEN_4940;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2b0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_688 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2b0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_688 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_688 <= _GEN_4941;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2b1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_689 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2b1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_689 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_689 <= _GEN_4942;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2b2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_690 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2b2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_690 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_690 <= _GEN_4943;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2b3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_691 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2b3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_691 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_691 <= _GEN_4944;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2b4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_692 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2b4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_692 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_692 <= _GEN_4945;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2b5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_693 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2b5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_693 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_693 <= _GEN_4946;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2b6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_694 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2b6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_694 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_694 <= _GEN_4947;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2b7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_695 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2b7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_695 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_695 <= _GEN_4948;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2b8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_696 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2b8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_696 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_696 <= _GEN_4949;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2b9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_697 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2b9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_697 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_697 <= _GEN_4950;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ba == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_698 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ba == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_698 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_698 <= _GEN_4951;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2bb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_699 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2bb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_699 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_699 <= _GEN_4952;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2bc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_700 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2bc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_700 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_700 <= _GEN_4953;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2bd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_701 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2bd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_701 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_701 <= _GEN_4954;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2be == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_702 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2be == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_702 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_702 <= _GEN_4955;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2bf == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_703 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2bf == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_703 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_703 <= _GEN_4956;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2c0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_704 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2c0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_704 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_704 <= _GEN_4957;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2c1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_705 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2c1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_705 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_705 <= _GEN_4958;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2c2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_706 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2c2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_706 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_706 <= _GEN_4959;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2c3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_707 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2c3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_707 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_707 <= _GEN_4960;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2c4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_708 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2c4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_708 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_708 <= _GEN_4961;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2c5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_709 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2c5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_709 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_709 <= _GEN_4962;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2c6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_710 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2c6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_710 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_710 <= _GEN_4963;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2c7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_711 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2c7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_711 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_711 <= _GEN_4964;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2c8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_712 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2c8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_712 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_712 <= _GEN_4965;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2c9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_713 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2c9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_713 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_713 <= _GEN_4966;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ca == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_714 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ca == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_714 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_714 <= _GEN_4967;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2cb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_715 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2cb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_715 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_715 <= _GEN_4968;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2cc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_716 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2cc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_716 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_716 <= _GEN_4969;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2cd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_717 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2cd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_717 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_717 <= _GEN_4970;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ce == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_718 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ce == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_718 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_718 <= _GEN_4971;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2cf == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_719 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2cf == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_719 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_719 <= _GEN_4972;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2d0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_720 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2d0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_720 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_720 <= _GEN_4973;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2d1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_721 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2d1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_721 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_721 <= _GEN_4974;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2d2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_722 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2d2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_722 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_722 <= _GEN_4975;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2d3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_723 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2d3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_723 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_723 <= _GEN_4976;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2d4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_724 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2d4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_724 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_724 <= _GEN_4977;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2d5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_725 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2d5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_725 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_725 <= _GEN_4978;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2d6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_726 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2d6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_726 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_726 <= _GEN_4979;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2d7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_727 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2d7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_727 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_727 <= _GEN_4980;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2d8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_728 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2d8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_728 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_728 <= _GEN_4981;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2d9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_729 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2d9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_729 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_729 <= _GEN_4982;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2da == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_730 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2da == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_730 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_730 <= _GEN_4983;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2db == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_731 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2db == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_731 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_731 <= _GEN_4984;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2dc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_732 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2dc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_732 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_732 <= _GEN_4985;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2dd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_733 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2dd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_733 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_733 <= _GEN_4986;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2de == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_734 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2de == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_734 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_734 <= _GEN_4987;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2df == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_735 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2df == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_735 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_735 <= _GEN_4988;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2e0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_736 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2e0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_736 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_736 <= _GEN_4989;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2e1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_737 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2e1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_737 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_737 <= _GEN_4990;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2e2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_738 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2e2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_738 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_738 <= _GEN_4991;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2e3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_739 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2e3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_739 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_739 <= _GEN_4992;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2e4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_740 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2e4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_740 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_740 <= _GEN_4993;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2e5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_741 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2e5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_741 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_741 <= _GEN_4994;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2e6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_742 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2e6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_742 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_742 <= _GEN_4995;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2e7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_743 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2e7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_743 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_743 <= _GEN_4996;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2e8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_744 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2e8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_744 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_744 <= _GEN_4997;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2e9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_745 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2e9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_745 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_745 <= _GEN_4998;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ea == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_746 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ea == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_746 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_746 <= _GEN_4999;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2eb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_747 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2eb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_747 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_747 <= _GEN_5000;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ec == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_748 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ec == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_748 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_748 <= _GEN_5001;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ed == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_749 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ed == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_749 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_749 <= _GEN_5002;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ee == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_750 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ee == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_750 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_750 <= _GEN_5003;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ef == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_751 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ef == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_751 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_751 <= _GEN_5004;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2f0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_752 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2f0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_752 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_752 <= _GEN_5005;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2f1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_753 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2f1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_753 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_753 <= _GEN_5006;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2f2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_754 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2f2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_754 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_754 <= _GEN_5007;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2f3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_755 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2f3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_755 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_755 <= _GEN_5008;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2f4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_756 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2f4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_756 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_756 <= _GEN_5009;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2f5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_757 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2f5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_757 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_757 <= _GEN_5010;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2f6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_758 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2f6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_758 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_758 <= _GEN_5011;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2f7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_759 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2f7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_759 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_759 <= _GEN_5012;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2f8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_760 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2f8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_760 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_760 <= _GEN_5013;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2f9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_761 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2f9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_761 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_761 <= _GEN_5014;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2fa == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_762 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2fa == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_762 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_762 <= _GEN_5015;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2fb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_763 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2fb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_763 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_763 <= _GEN_5016;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2fc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_764 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2fc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_764 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_764 <= _GEN_5017;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2fd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_765 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2fd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_765 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_765 <= _GEN_5018;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2fe == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_766 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2fe == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_766 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_766 <= _GEN_5019;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h2ff == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_767 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h2ff == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_767 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_767 <= _GEN_5020;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h300 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_768 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h300 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_768 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_768 <= _GEN_5021;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h301 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_769 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h301 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_769 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_769 <= _GEN_5022;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h302 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_770 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h302 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_770 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_770 <= _GEN_5023;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h303 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_771 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h303 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_771 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_771 <= _GEN_5024;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h304 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_772 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h304 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_772 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_772 <= _GEN_5025;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h305 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_773 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h305 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_773 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_773 <= _GEN_5026;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h306 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_774 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h306 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_774 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_774 <= _GEN_5027;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h307 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_775 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h307 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_775 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_775 <= _GEN_5028;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h308 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_776 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h308 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_776 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_776 <= _GEN_5029;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h309 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_777 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h309 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_777 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_777 <= _GEN_5030;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h30a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_778 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h30a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_778 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_778 <= _GEN_5031;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h30b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_779 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h30b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_779 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_779 <= _GEN_5032;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h30c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_780 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h30c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_780 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_780 <= _GEN_5033;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h30d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_781 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h30d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_781 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_781 <= _GEN_5034;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h30e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_782 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h30e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_782 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_782 <= _GEN_5035;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h30f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_783 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h30f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_783 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_783 <= _GEN_5036;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h310 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_784 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h310 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_784 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_784 <= _GEN_5037;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h311 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_785 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h311 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_785 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_785 <= _GEN_5038;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h312 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_786 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h312 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_786 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_786 <= _GEN_5039;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h313 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_787 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h313 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_787 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_787 <= _GEN_5040;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h314 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_788 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h314 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_788 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_788 <= _GEN_5041;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h315 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_789 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h315 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_789 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_789 <= _GEN_5042;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h316 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_790 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h316 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_790 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_790 <= _GEN_5043;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h317 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_791 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h317 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_791 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_791 <= _GEN_5044;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h318 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_792 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h318 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_792 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_792 <= _GEN_5045;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h319 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_793 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h319 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_793 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_793 <= _GEN_5046;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h31a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_794 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h31a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_794 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_794 <= _GEN_5047;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h31b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_795 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h31b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_795 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_795 <= _GEN_5048;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h31c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_796 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h31c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_796 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_796 <= _GEN_5049;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h31d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_797 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h31d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_797 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_797 <= _GEN_5050;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h31e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_798 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h31e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_798 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_798 <= _GEN_5051;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h31f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_799 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h31f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_799 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_799 <= _GEN_5052;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h320 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_800 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h320 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_800 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_800 <= _GEN_5053;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h321 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_801 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h321 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_801 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_801 <= _GEN_5054;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h322 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_802 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h322 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_802 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_802 <= _GEN_5055;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h323 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_803 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h323 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_803 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_803 <= _GEN_5056;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h324 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_804 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h324 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_804 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_804 <= _GEN_5057;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h325 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_805 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h325 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_805 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_805 <= _GEN_5058;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h326 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_806 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h326 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_806 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_806 <= _GEN_5059;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h327 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_807 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h327 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_807 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_807 <= _GEN_5060;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h328 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_808 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h328 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_808 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_808 <= _GEN_5061;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h329 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_809 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h329 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_809 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_809 <= _GEN_5062;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h32a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_810 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h32a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_810 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_810 <= _GEN_5063;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h32b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_811 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h32b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_811 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_811 <= _GEN_5064;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h32c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_812 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h32c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_812 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_812 <= _GEN_5065;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h32d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_813 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h32d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_813 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_813 <= _GEN_5066;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h32e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_814 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h32e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_814 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_814 <= _GEN_5067;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h32f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_815 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h32f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_815 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_815 <= _GEN_5068;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h330 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_816 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h330 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_816 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_816 <= _GEN_5069;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h331 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_817 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h331 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_817 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_817 <= _GEN_5070;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h332 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_818 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h332 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_818 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_818 <= _GEN_5071;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h333 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_819 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h333 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_819 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_819 <= _GEN_5072;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h334 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_820 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h334 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_820 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_820 <= _GEN_5073;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h335 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_821 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h335 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_821 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_821 <= _GEN_5074;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h336 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_822 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h336 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_822 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_822 <= _GEN_5075;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h337 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_823 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h337 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_823 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_823 <= _GEN_5076;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h338 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_824 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h338 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_824 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_824 <= _GEN_5077;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h339 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_825 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h339 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_825 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_825 <= _GEN_5078;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h33a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_826 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h33a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_826 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_826 <= _GEN_5079;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h33b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_827 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h33b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_827 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_827 <= _GEN_5080;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h33c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_828 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h33c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_828 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_828 <= _GEN_5081;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h33d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_829 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h33d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_829 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_829 <= _GEN_5082;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h33e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_830 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h33e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_830 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_830 <= _GEN_5083;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h33f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_831 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h33f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_831 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_831 <= _GEN_5084;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h340 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_832 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h340 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_832 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_832 <= _GEN_5085;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h341 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_833 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h341 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_833 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_833 <= _GEN_5086;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h342 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_834 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h342 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_834 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_834 <= _GEN_5087;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h343 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_835 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h343 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_835 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_835 <= _GEN_5088;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h344 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_836 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h344 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_836 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_836 <= _GEN_5089;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h345 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_837 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h345 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_837 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_837 <= _GEN_5090;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h346 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_838 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h346 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_838 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_838 <= _GEN_5091;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h347 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_839 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h347 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_839 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_839 <= _GEN_5092;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h348 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_840 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h348 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_840 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_840 <= _GEN_5093;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h349 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_841 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h349 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_841 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_841 <= _GEN_5094;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h34a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_842 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h34a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_842 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_842 <= _GEN_5095;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h34b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_843 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h34b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_843 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_843 <= _GEN_5096;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h34c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_844 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h34c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_844 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_844 <= _GEN_5097;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h34d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_845 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h34d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_845 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_845 <= _GEN_5098;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h34e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_846 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h34e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_846 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_846 <= _GEN_5099;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h34f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_847 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h34f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_847 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_847 <= _GEN_5100;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h350 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_848 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h350 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_848 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_848 <= _GEN_5101;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h351 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_849 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h351 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_849 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_849 <= _GEN_5102;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h352 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_850 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h352 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_850 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_850 <= _GEN_5103;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h353 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_851 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h353 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_851 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_851 <= _GEN_5104;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h354 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_852 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h354 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_852 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_852 <= _GEN_5105;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h355 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_853 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h355 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_853 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_853 <= _GEN_5106;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h356 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_854 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h356 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_854 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_854 <= _GEN_5107;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h357 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_855 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h357 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_855 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_855 <= _GEN_5108;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h358 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_856 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h358 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_856 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_856 <= _GEN_5109;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h359 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_857 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h359 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_857 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_857 <= _GEN_5110;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h35a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_858 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h35a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_858 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_858 <= _GEN_5111;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h35b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_859 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h35b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_859 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_859 <= _GEN_5112;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h35c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_860 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h35c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_860 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_860 <= _GEN_5113;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h35d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_861 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h35d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_861 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_861 <= _GEN_5114;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h35e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_862 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h35e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_862 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_862 <= _GEN_5115;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h35f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_863 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h35f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_863 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_863 <= _GEN_5116;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h360 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_864 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h360 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_864 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_864 <= _GEN_5117;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h361 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_865 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h361 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_865 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_865 <= _GEN_5118;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h362 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_866 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h362 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_866 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_866 <= _GEN_5119;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h363 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_867 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h363 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_867 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_867 <= _GEN_5120;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h364 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_868 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h364 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_868 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_868 <= _GEN_5121;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h365 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_869 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h365 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_869 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_869 <= _GEN_5122;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h366 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_870 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h366 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_870 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_870 <= _GEN_5123;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h367 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_871 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h367 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_871 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_871 <= _GEN_5124;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h368 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_872 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h368 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_872 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_872 <= _GEN_5125;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h369 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_873 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h369 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_873 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_873 <= _GEN_5126;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h36a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_874 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h36a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_874 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_874 <= _GEN_5127;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h36b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_875 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h36b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_875 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_875 <= _GEN_5128;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h36c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_876 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h36c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_876 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_876 <= _GEN_5129;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h36d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_877 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h36d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_877 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_877 <= _GEN_5130;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h36e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_878 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h36e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_878 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_878 <= _GEN_5131;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h36f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_879 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h36f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_879 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_879 <= _GEN_5132;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h370 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_880 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h370 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_880 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_880 <= _GEN_5133;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h371 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_881 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h371 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_881 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_881 <= _GEN_5134;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h372 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_882 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h372 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_882 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_882 <= _GEN_5135;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h373 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_883 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h373 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_883 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_883 <= _GEN_5136;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h374 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_884 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h374 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_884 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_884 <= _GEN_5137;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h375 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_885 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h375 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_885 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_885 <= _GEN_5138;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h376 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_886 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h376 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_886 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_886 <= _GEN_5139;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h377 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_887 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h377 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_887 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_887 <= _GEN_5140;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h378 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_888 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h378 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_888 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_888 <= _GEN_5141;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h379 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_889 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h379 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_889 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_889 <= _GEN_5142;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h37a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_890 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h37a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_890 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_890 <= _GEN_5143;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h37b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_891 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h37b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_891 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_891 <= _GEN_5144;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h37c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_892 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h37c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_892 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_892 <= _GEN_5145;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h37d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_893 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h37d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_893 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_893 <= _GEN_5146;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h37e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_894 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h37e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_894 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_894 <= _GEN_5147;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h37f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_895 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h37f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_895 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_895 <= _GEN_5148;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h380 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_896 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h380 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_896 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_896 <= _GEN_5149;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h381 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_897 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h381 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_897 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_897 <= _GEN_5150;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h382 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_898 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h382 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_898 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_898 <= _GEN_5151;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h383 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_899 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h383 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_899 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_899 <= _GEN_5152;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h384 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_900 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h384 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_900 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_900 <= _GEN_5153;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h385 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_901 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h385 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_901 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_901 <= _GEN_5154;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h386 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_902 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h386 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_902 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_902 <= _GEN_5155;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h387 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_903 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h387 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_903 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_903 <= _GEN_5156;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h388 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_904 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h388 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_904 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_904 <= _GEN_5157;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h389 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_905 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h389 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_905 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_905 <= _GEN_5158;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h38a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_906 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h38a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_906 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_906 <= _GEN_5159;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h38b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_907 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h38b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_907 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_907 <= _GEN_5160;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h38c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_908 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h38c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_908 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_908 <= _GEN_5161;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h38d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_909 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h38d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_909 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_909 <= _GEN_5162;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h38e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_910 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h38e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_910 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_910 <= _GEN_5163;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h38f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_911 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h38f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_911 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_911 <= _GEN_5164;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h390 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_912 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h390 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_912 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_912 <= _GEN_5165;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h391 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_913 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h391 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_913 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_913 <= _GEN_5166;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h392 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_914 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h392 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_914 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_914 <= _GEN_5167;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h393 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_915 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h393 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_915 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_915 <= _GEN_5168;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h394 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_916 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h394 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_916 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_916 <= _GEN_5169;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h395 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_917 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h395 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_917 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_917 <= _GEN_5170;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h396 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_918 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h396 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_918 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_918 <= _GEN_5171;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h397 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_919 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h397 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_919 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_919 <= _GEN_5172;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h398 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_920 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h398 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_920 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_920 <= _GEN_5173;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h399 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_921 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h399 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_921 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_921 <= _GEN_5174;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h39a == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_922 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h39a == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_922 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_922 <= _GEN_5175;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h39b == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_923 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h39b == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_923 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_923 <= _GEN_5176;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h39c == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_924 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h39c == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_924 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_924 <= _GEN_5177;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h39d == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_925 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h39d == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_925 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_925 <= _GEN_5178;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h39e == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_926 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h39e == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_926 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_926 <= _GEN_5179;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h39f == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_927 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h39f == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_927 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_927 <= _GEN_5180;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3a0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_928 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3a0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_928 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_928 <= _GEN_5181;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3a1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_929 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3a1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_929 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_929 <= _GEN_5182;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3a2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_930 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3a2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_930 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_930 <= _GEN_5183;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3a3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_931 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3a3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_931 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_931 <= _GEN_5184;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3a4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_932 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3a4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_932 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_932 <= _GEN_5185;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3a5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_933 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3a5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_933 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_933 <= _GEN_5186;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3a6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_934 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3a6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_934 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_934 <= _GEN_5187;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3a7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_935 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3a7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_935 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_935 <= _GEN_5188;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3a8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_936 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3a8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_936 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_936 <= _GEN_5189;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3a9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_937 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3a9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_937 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_937 <= _GEN_5190;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3aa == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_938 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3aa == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_938 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_938 <= _GEN_5191;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ab == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_939 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ab == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_939 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_939 <= _GEN_5192;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ac == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_940 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ac == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_940 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_940 <= _GEN_5193;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ad == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_941 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ad == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_941 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_941 <= _GEN_5194;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ae == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_942 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ae == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_942 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_942 <= _GEN_5195;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3af == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_943 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3af == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_943 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_943 <= _GEN_5196;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3b0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_944 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3b0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_944 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_944 <= _GEN_5197;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3b1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_945 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3b1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_945 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_945 <= _GEN_5198;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3b2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_946 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3b2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_946 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_946 <= _GEN_5199;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3b3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_947 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3b3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_947 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_947 <= _GEN_5200;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3b4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_948 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3b4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_948 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_948 <= _GEN_5201;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3b5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_949 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3b5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_949 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_949 <= _GEN_5202;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3b6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_950 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3b6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_950 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_950 <= _GEN_5203;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3b7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_951 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3b7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_951 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_951 <= _GEN_5204;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3b8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_952 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3b8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_952 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_952 <= _GEN_5205;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3b9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_953 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3b9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_953 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_953 <= _GEN_5206;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ba == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_954 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ba == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_954 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_954 <= _GEN_5207;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3bb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_955 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3bb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_955 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_955 <= _GEN_5208;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3bc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_956 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3bc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_956 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_956 <= _GEN_5209;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3bd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_957 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3bd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_957 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_957 <= _GEN_5210;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3be == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_958 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3be == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_958 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_958 <= _GEN_5211;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3bf == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_959 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3bf == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_959 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_959 <= _GEN_5212;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3c0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_960 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3c0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_960 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_960 <= _GEN_5213;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3c1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_961 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3c1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_961 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_961 <= _GEN_5214;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3c2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_962 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3c2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_962 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_962 <= _GEN_5215;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3c3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_963 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3c3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_963 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_963 <= _GEN_5216;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3c4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_964 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3c4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_964 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_964 <= _GEN_5217;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3c5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_965 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3c5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_965 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_965 <= _GEN_5218;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3c6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_966 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3c6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_966 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_966 <= _GEN_5219;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3c7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_967 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3c7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_967 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_967 <= _GEN_5220;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3c8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_968 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3c8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_968 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_968 <= _GEN_5221;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3c9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_969 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3c9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_969 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_969 <= _GEN_5222;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ca == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_970 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ca == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_970 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_970 <= _GEN_5223;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3cb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_971 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3cb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_971 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_971 <= _GEN_5224;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3cc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_972 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3cc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_972 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_972 <= _GEN_5225;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3cd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_973 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3cd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_973 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_973 <= _GEN_5226;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ce == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_974 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ce == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_974 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_974 <= _GEN_5227;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3cf == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_975 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3cf == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_975 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_975 <= _GEN_5228;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3d0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_976 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3d0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_976 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_976 <= _GEN_5229;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3d1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_977 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3d1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_977 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_977 <= _GEN_5230;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3d2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_978 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3d2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_978 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_978 <= _GEN_5231;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3d3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_979 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3d3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_979 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_979 <= _GEN_5232;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3d4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_980 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3d4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_980 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_980 <= _GEN_5233;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3d5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_981 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3d5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_981 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_981 <= _GEN_5234;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3d6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_982 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3d6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_982 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_982 <= _GEN_5235;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3d7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_983 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3d7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_983 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_983 <= _GEN_5236;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3d8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_984 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3d8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_984 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_984 <= _GEN_5237;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3d9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_985 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3d9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_985 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_985 <= _GEN_5238;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3da == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_986 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3da == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_986 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_986 <= _GEN_5239;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3db == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_987 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3db == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_987 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_987 <= _GEN_5240;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3dc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_988 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3dc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_988 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_988 <= _GEN_5241;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3dd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_989 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3dd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_989 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_989 <= _GEN_5242;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3de == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_990 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3de == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_990 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_990 <= _GEN_5243;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3df == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_991 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3df == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_991 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_991 <= _GEN_5244;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3e0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_992 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3e0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_992 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_992 <= _GEN_5245;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3e1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_993 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3e1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_993 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_993 <= _GEN_5246;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3e2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_994 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3e2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_994 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_994 <= _GEN_5247;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3e3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_995 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3e3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_995 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_995 <= _GEN_5248;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3e4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_996 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3e4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_996 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_996 <= _GEN_5249;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3e5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_997 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3e5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_997 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_997 <= _GEN_5250;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3e6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_998 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3e6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_998 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_998 <= _GEN_5251;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3e7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_999 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3e7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_999 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_999 <= _GEN_5252;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3e8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1000 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3e8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1000 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1000 <= _GEN_5253;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3e9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1001 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3e9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1001 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1001 <= _GEN_5254;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ea == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1002 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ea == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1002 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1002 <= _GEN_5255;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3eb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1003 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3eb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1003 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1003 <= _GEN_5256;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ec == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1004 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ec == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1004 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1004 <= _GEN_5257;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ed == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1005 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ed == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1005 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1005 <= _GEN_5258;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ee == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1006 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ee == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1006 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1006 <= _GEN_5259;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ef == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1007 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ef == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1007 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1007 <= _GEN_5260;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3f0 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1008 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3f0 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1008 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1008 <= _GEN_5261;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3f1 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1009 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3f1 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1009 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1009 <= _GEN_5262;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3f2 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1010 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3f2 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1010 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1010 <= _GEN_5263;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3f3 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1011 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3f3 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1011 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1011 <= _GEN_5264;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3f4 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1012 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3f4 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1012 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1012 <= _GEN_5265;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3f5 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1013 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3f5 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1013 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1013 <= _GEN_5266;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3f6 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1014 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3f6 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1014 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1014 <= _GEN_5267;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3f7 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1015 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3f7 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1015 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1015 <= _GEN_5268;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3f8 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1016 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3f8 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1016 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1016 <= _GEN_5269;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3f9 == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1017 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3f9 == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1017 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1017 <= _GEN_5270;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3fa == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1018 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3fa == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1018 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1018 <= _GEN_5271;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3fb == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1019 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3fb == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1019 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1019 <= _GEN_5272;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3fc == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1020 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3fc == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1020 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1020 <= _GEN_5273;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3fd == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1021 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3fd == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1021 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1021 <= _GEN_5274;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3fe == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1022 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3fe == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1022 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1022 <= _GEN_5275;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      if (10'h3ff == io_rvfi_mem_addr_in_1) begin // @[CPU.scala 75:39]
        DMemory_1023 <= io_rvfi_mem_data_in_1; // @[CPU.scala 75:39]
      end else if (10'h3ff == io_rvfi_mem_addr_in_0) begin // @[CPU.scala 75:39]
        DMemory_1023 <= io_rvfi_mem_data_in_0; // @[CPU.scala 75:39]
      end
    end else if (!(_bypassAFromMEM_T_3)) begin // @[CPU.scala 200:29]
      if (!(_stall_T)) begin // @[CPU.scala 202:32]
        if (EXMEMop == 7'h23) begin // @[CPU.scala 204:32]
          DMemory_1023 <= _GEN_5276;
        end
      end
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      IMemory_0 <= io_rvfi_insn_in_0; // @[CPU.scala 72:18]
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      IMemory_1 <= io_rvfi_insn_in_1; // @[CPU.scala 72:18]
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      IMemory_2 <= io_rvfi_insn_in_2; // @[CPU.scala 72:18]
    end
    if (io_rvfi_rst) begin // @[CPU.scala 61:21]
      IMemory_3 <= io_rvfi_insn_in_3; // @[CPU.scala 72:18]
    end
    if (reset) begin // @[CPU.scala 54:49]
      IFIDIR <= 32'h13; // @[CPU.scala 54:49]
    end else if (!(io_rvfi_rst)) begin // @[CPU.scala 61:21]
      if (~stall) begin // @[CPU.scala 121:27]
        if (~takeBranch) begin // @[CPU.scala 122:34]
          IFIDIR <= _GEN_3135; // @[CPU.scala 125:16]
        end else begin
          IFIDIR <= 32'h13; // @[CPU.scala 129:16]
        end
      end
    end
    if (reset) begin // @[CPU.scala 54:49]
      IDEXIR <= 32'h13; // @[CPU.scala 54:49]
    end else if (!(io_rvfi_rst)) begin // @[CPU.scala 61:21]
      if (~stall) begin // @[CPU.scala 121:27]
        IDEXIR <= IFIDIR; // @[CPU.scala 174:14]
      end else begin
        IDEXIR <= 32'h13; // @[CPU.scala 176:14]
      end
    end
    if (reset) begin // @[CPU.scala 54:49]
      EXMEMIR <= 32'h13; // @[CPU.scala 54:49]
    end else if (!(io_rvfi_rst)) begin // @[CPU.scala 61:21]
      EXMEMIR <= IDEXIR; // @[CPU.scala 196:13]
    end
    if (reset) begin // @[CPU.scala 54:49]
      MEMWBIR <= 32'h13; // @[CPU.scala 54:49]
    end else if (!(io_rvfi_rst)) begin // @[CPU.scala 61:21]
      MEMWBIR <= EXMEMIR; // @[CPU.scala 208:13]
    end
    if (reset) begin // @[CPU.scala 57:22]
      CurPC <= 64'h0; // @[CPU.scala 57:22]
    end else if (!(io_rvfi_rst)) begin // @[CPU.scala 61:21]
      if (~stall) begin // @[CPU.scala 121:27]
        CurPC <= PC; // @[CPU.scala 145:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  PC = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  Regs_0 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  Regs_1 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  Regs_2 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  Regs_3 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  Regs_4 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  Regs_5 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  Regs_6 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  Regs_7 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  Regs_8 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  Regs_9 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  Regs_10 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  Regs_11 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  Regs_12 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  Regs_13 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  Regs_14 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  Regs_15 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  Regs_16 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  Regs_17 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  Regs_18 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  Regs_19 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  Regs_20 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  Regs_21 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  Regs_22 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  Regs_23 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  Regs_24 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  Regs_25 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  Regs_26 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  Regs_27 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  Regs_28 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  Regs_29 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  Regs_30 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  Regs_31 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  IDEXA = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  IDEXB = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  EXMEMB = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  EXMEMALUOut = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  MEMWBValue = _RAND_37[63:0];
  _RAND_38 = {1{`RANDOM}};
  DMemory_0 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  DMemory_1 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  DMemory_2 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  DMemory_3 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  DMemory_4 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  DMemory_5 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  DMemory_6 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  DMemory_7 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  DMemory_8 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  DMemory_9 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  DMemory_10 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  DMemory_11 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  DMemory_12 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  DMemory_13 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  DMemory_14 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  DMemory_15 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  DMemory_16 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  DMemory_17 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  DMemory_18 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  DMemory_19 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  DMemory_20 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  DMemory_21 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  DMemory_22 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  DMemory_23 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  DMemory_24 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  DMemory_25 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  DMemory_26 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  DMemory_27 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  DMemory_28 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  DMemory_29 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  DMemory_30 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  DMemory_31 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  DMemory_32 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  DMemory_33 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  DMemory_34 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  DMemory_35 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  DMemory_36 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  DMemory_37 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  DMemory_38 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  DMemory_39 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  DMemory_40 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  DMemory_41 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  DMemory_42 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  DMemory_43 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  DMemory_44 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  DMemory_45 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  DMemory_46 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  DMemory_47 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  DMemory_48 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  DMemory_49 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  DMemory_50 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  DMemory_51 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  DMemory_52 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  DMemory_53 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  DMemory_54 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  DMemory_55 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  DMemory_56 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  DMemory_57 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  DMemory_58 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  DMemory_59 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  DMemory_60 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  DMemory_61 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  DMemory_62 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  DMemory_63 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  DMemory_64 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  DMemory_65 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  DMemory_66 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  DMemory_67 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  DMemory_68 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  DMemory_69 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  DMemory_70 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  DMemory_71 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  DMemory_72 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  DMemory_73 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  DMemory_74 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  DMemory_75 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  DMemory_76 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  DMemory_77 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  DMemory_78 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  DMemory_79 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  DMemory_80 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  DMemory_81 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  DMemory_82 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  DMemory_83 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  DMemory_84 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  DMemory_85 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  DMemory_86 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  DMemory_87 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  DMemory_88 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  DMemory_89 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  DMemory_90 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  DMemory_91 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  DMemory_92 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  DMemory_93 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  DMemory_94 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  DMemory_95 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  DMemory_96 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  DMemory_97 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  DMemory_98 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  DMemory_99 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  DMemory_100 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  DMemory_101 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  DMemory_102 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  DMemory_103 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  DMemory_104 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  DMemory_105 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  DMemory_106 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  DMemory_107 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  DMemory_108 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  DMemory_109 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  DMemory_110 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  DMemory_111 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  DMemory_112 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  DMemory_113 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  DMemory_114 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  DMemory_115 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  DMemory_116 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  DMemory_117 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  DMemory_118 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  DMemory_119 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  DMemory_120 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  DMemory_121 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  DMemory_122 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  DMemory_123 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  DMemory_124 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  DMemory_125 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  DMemory_126 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  DMemory_127 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  DMemory_128 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  DMemory_129 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  DMemory_130 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  DMemory_131 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  DMemory_132 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  DMemory_133 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  DMemory_134 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  DMemory_135 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  DMemory_136 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  DMemory_137 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  DMemory_138 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  DMemory_139 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  DMemory_140 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  DMemory_141 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  DMemory_142 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  DMemory_143 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  DMemory_144 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  DMemory_145 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  DMemory_146 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  DMemory_147 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  DMemory_148 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  DMemory_149 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  DMemory_150 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  DMemory_151 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  DMemory_152 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  DMemory_153 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  DMemory_154 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  DMemory_155 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  DMemory_156 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  DMemory_157 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  DMemory_158 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  DMemory_159 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  DMemory_160 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  DMemory_161 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  DMemory_162 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  DMemory_163 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  DMemory_164 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  DMemory_165 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  DMemory_166 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  DMemory_167 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  DMemory_168 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  DMemory_169 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  DMemory_170 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  DMemory_171 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  DMemory_172 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  DMemory_173 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  DMemory_174 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  DMemory_175 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  DMemory_176 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  DMemory_177 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  DMemory_178 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  DMemory_179 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  DMemory_180 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  DMemory_181 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  DMemory_182 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  DMemory_183 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  DMemory_184 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  DMemory_185 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  DMemory_186 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  DMemory_187 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  DMemory_188 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  DMemory_189 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  DMemory_190 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  DMemory_191 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  DMemory_192 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  DMemory_193 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  DMemory_194 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  DMemory_195 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  DMemory_196 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  DMemory_197 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  DMemory_198 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  DMemory_199 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  DMemory_200 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  DMemory_201 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  DMemory_202 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  DMemory_203 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  DMemory_204 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  DMemory_205 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  DMemory_206 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  DMemory_207 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  DMemory_208 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  DMemory_209 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  DMemory_210 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  DMemory_211 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  DMemory_212 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  DMemory_213 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  DMemory_214 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  DMemory_215 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  DMemory_216 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  DMemory_217 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  DMemory_218 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  DMemory_219 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  DMemory_220 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  DMemory_221 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  DMemory_222 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  DMemory_223 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  DMemory_224 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  DMemory_225 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  DMemory_226 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  DMemory_227 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  DMemory_228 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  DMemory_229 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  DMemory_230 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  DMemory_231 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  DMemory_232 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  DMemory_233 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  DMemory_234 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  DMemory_235 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  DMemory_236 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  DMemory_237 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  DMemory_238 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  DMemory_239 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  DMemory_240 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  DMemory_241 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  DMemory_242 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  DMemory_243 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  DMemory_244 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  DMemory_245 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  DMemory_246 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  DMemory_247 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  DMemory_248 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  DMemory_249 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  DMemory_250 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  DMemory_251 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  DMemory_252 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  DMemory_253 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  DMemory_254 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  DMemory_255 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  DMemory_256 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  DMemory_257 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  DMemory_258 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  DMemory_259 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  DMemory_260 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  DMemory_261 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  DMemory_262 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  DMemory_263 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  DMemory_264 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  DMemory_265 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  DMemory_266 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  DMemory_267 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  DMemory_268 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  DMemory_269 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  DMemory_270 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  DMemory_271 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  DMemory_272 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  DMemory_273 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  DMemory_274 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  DMemory_275 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  DMemory_276 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  DMemory_277 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  DMemory_278 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  DMemory_279 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  DMemory_280 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  DMemory_281 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  DMemory_282 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  DMemory_283 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  DMemory_284 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  DMemory_285 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  DMemory_286 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  DMemory_287 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  DMemory_288 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  DMemory_289 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  DMemory_290 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  DMemory_291 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  DMemory_292 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  DMemory_293 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  DMemory_294 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  DMemory_295 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  DMemory_296 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  DMemory_297 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  DMemory_298 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  DMemory_299 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  DMemory_300 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  DMemory_301 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  DMemory_302 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  DMemory_303 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  DMemory_304 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  DMemory_305 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  DMemory_306 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  DMemory_307 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  DMemory_308 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  DMemory_309 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  DMemory_310 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  DMemory_311 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  DMemory_312 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  DMemory_313 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  DMemory_314 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  DMemory_315 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  DMemory_316 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  DMemory_317 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  DMemory_318 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  DMemory_319 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  DMemory_320 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  DMemory_321 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  DMemory_322 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  DMemory_323 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  DMemory_324 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  DMemory_325 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  DMemory_326 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  DMemory_327 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  DMemory_328 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  DMemory_329 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  DMemory_330 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  DMemory_331 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  DMemory_332 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  DMemory_333 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  DMemory_334 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  DMemory_335 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  DMemory_336 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  DMemory_337 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  DMemory_338 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  DMemory_339 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  DMemory_340 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  DMemory_341 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  DMemory_342 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  DMemory_343 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  DMemory_344 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  DMemory_345 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  DMemory_346 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  DMemory_347 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  DMemory_348 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  DMemory_349 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  DMemory_350 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  DMemory_351 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  DMemory_352 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  DMemory_353 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  DMemory_354 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  DMemory_355 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  DMemory_356 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  DMemory_357 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  DMemory_358 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  DMemory_359 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  DMemory_360 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  DMemory_361 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  DMemory_362 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  DMemory_363 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  DMemory_364 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  DMemory_365 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  DMemory_366 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  DMemory_367 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  DMemory_368 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  DMemory_369 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  DMemory_370 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  DMemory_371 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  DMemory_372 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  DMemory_373 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  DMemory_374 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  DMemory_375 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  DMemory_376 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  DMemory_377 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  DMemory_378 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  DMemory_379 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  DMemory_380 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  DMemory_381 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  DMemory_382 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  DMemory_383 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  DMemory_384 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  DMemory_385 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  DMemory_386 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  DMemory_387 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  DMemory_388 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  DMemory_389 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  DMemory_390 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  DMemory_391 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  DMemory_392 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  DMemory_393 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  DMemory_394 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  DMemory_395 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  DMemory_396 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  DMemory_397 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  DMemory_398 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  DMemory_399 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  DMemory_400 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  DMemory_401 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  DMemory_402 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  DMemory_403 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  DMemory_404 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  DMemory_405 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  DMemory_406 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  DMemory_407 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  DMemory_408 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  DMemory_409 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  DMemory_410 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  DMemory_411 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  DMemory_412 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  DMemory_413 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  DMemory_414 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  DMemory_415 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  DMemory_416 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  DMemory_417 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  DMemory_418 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  DMemory_419 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  DMemory_420 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  DMemory_421 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  DMemory_422 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  DMemory_423 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  DMemory_424 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  DMemory_425 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  DMemory_426 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  DMemory_427 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  DMemory_428 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  DMemory_429 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  DMemory_430 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  DMemory_431 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  DMemory_432 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  DMemory_433 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  DMemory_434 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  DMemory_435 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  DMemory_436 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  DMemory_437 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  DMemory_438 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  DMemory_439 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  DMemory_440 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  DMemory_441 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  DMemory_442 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  DMemory_443 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  DMemory_444 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  DMemory_445 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  DMemory_446 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  DMemory_447 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  DMemory_448 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  DMemory_449 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  DMemory_450 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  DMemory_451 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  DMemory_452 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  DMemory_453 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  DMemory_454 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  DMemory_455 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  DMemory_456 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  DMemory_457 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  DMemory_458 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  DMemory_459 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  DMemory_460 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  DMemory_461 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  DMemory_462 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  DMemory_463 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  DMemory_464 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  DMemory_465 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  DMemory_466 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  DMemory_467 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  DMemory_468 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  DMemory_469 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  DMemory_470 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  DMemory_471 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  DMemory_472 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  DMemory_473 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  DMemory_474 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  DMemory_475 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  DMemory_476 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  DMemory_477 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  DMemory_478 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  DMemory_479 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  DMemory_480 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  DMemory_481 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  DMemory_482 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  DMemory_483 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  DMemory_484 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  DMemory_485 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  DMemory_486 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  DMemory_487 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  DMemory_488 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  DMemory_489 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  DMemory_490 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  DMemory_491 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  DMemory_492 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  DMemory_493 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  DMemory_494 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  DMemory_495 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  DMemory_496 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  DMemory_497 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  DMemory_498 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  DMemory_499 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  DMemory_500 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  DMemory_501 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  DMemory_502 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  DMemory_503 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  DMemory_504 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  DMemory_505 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  DMemory_506 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  DMemory_507 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  DMemory_508 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  DMemory_509 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  DMemory_510 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  DMemory_511 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  DMemory_512 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  DMemory_513 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  DMemory_514 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  DMemory_515 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  DMemory_516 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  DMemory_517 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  DMemory_518 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  DMemory_519 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  DMemory_520 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  DMemory_521 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  DMemory_522 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  DMemory_523 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  DMemory_524 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  DMemory_525 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  DMemory_526 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  DMemory_527 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  DMemory_528 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  DMemory_529 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  DMemory_530 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  DMemory_531 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  DMemory_532 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  DMemory_533 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  DMemory_534 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  DMemory_535 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  DMemory_536 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  DMemory_537 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  DMemory_538 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  DMemory_539 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  DMemory_540 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  DMemory_541 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  DMemory_542 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  DMemory_543 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  DMemory_544 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  DMemory_545 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  DMemory_546 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  DMemory_547 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  DMemory_548 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  DMemory_549 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  DMemory_550 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  DMemory_551 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  DMemory_552 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  DMemory_553 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  DMemory_554 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  DMemory_555 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  DMemory_556 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  DMemory_557 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  DMemory_558 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  DMemory_559 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  DMemory_560 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  DMemory_561 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  DMemory_562 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  DMemory_563 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  DMemory_564 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  DMemory_565 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  DMemory_566 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  DMemory_567 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  DMemory_568 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  DMemory_569 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  DMemory_570 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  DMemory_571 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  DMemory_572 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  DMemory_573 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  DMemory_574 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  DMemory_575 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  DMemory_576 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  DMemory_577 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  DMemory_578 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  DMemory_579 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  DMemory_580 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  DMemory_581 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  DMemory_582 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  DMemory_583 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  DMemory_584 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  DMemory_585 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  DMemory_586 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  DMemory_587 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  DMemory_588 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  DMemory_589 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  DMemory_590 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  DMemory_591 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  DMemory_592 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  DMemory_593 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  DMemory_594 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  DMemory_595 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  DMemory_596 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  DMemory_597 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  DMemory_598 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  DMemory_599 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  DMemory_600 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  DMemory_601 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  DMemory_602 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  DMemory_603 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  DMemory_604 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  DMemory_605 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  DMemory_606 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  DMemory_607 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  DMemory_608 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  DMemory_609 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  DMemory_610 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  DMemory_611 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  DMemory_612 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  DMemory_613 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  DMemory_614 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  DMemory_615 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  DMemory_616 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  DMemory_617 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  DMemory_618 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  DMemory_619 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  DMemory_620 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  DMemory_621 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  DMemory_622 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  DMemory_623 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  DMemory_624 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  DMemory_625 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  DMemory_626 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  DMemory_627 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  DMemory_628 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  DMemory_629 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  DMemory_630 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  DMemory_631 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  DMemory_632 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  DMemory_633 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  DMemory_634 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  DMemory_635 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  DMemory_636 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  DMemory_637 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  DMemory_638 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  DMemory_639 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  DMemory_640 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  DMemory_641 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  DMemory_642 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  DMemory_643 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  DMemory_644 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  DMemory_645 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  DMemory_646 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  DMemory_647 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  DMemory_648 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  DMemory_649 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  DMemory_650 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  DMemory_651 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  DMemory_652 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  DMemory_653 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  DMemory_654 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  DMemory_655 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  DMemory_656 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  DMemory_657 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  DMemory_658 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  DMemory_659 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  DMemory_660 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  DMemory_661 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  DMemory_662 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  DMemory_663 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  DMemory_664 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  DMemory_665 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  DMemory_666 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  DMemory_667 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  DMemory_668 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  DMemory_669 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  DMemory_670 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  DMemory_671 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  DMemory_672 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  DMemory_673 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  DMemory_674 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  DMemory_675 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  DMemory_676 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  DMemory_677 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  DMemory_678 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  DMemory_679 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  DMemory_680 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  DMemory_681 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  DMemory_682 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  DMemory_683 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  DMemory_684 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  DMemory_685 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  DMemory_686 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  DMemory_687 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  DMemory_688 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  DMemory_689 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  DMemory_690 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  DMemory_691 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  DMemory_692 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  DMemory_693 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  DMemory_694 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  DMemory_695 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  DMemory_696 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  DMemory_697 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  DMemory_698 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  DMemory_699 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  DMemory_700 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  DMemory_701 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  DMemory_702 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  DMemory_703 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  DMemory_704 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  DMemory_705 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  DMemory_706 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  DMemory_707 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  DMemory_708 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  DMemory_709 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  DMemory_710 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  DMemory_711 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  DMemory_712 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  DMemory_713 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  DMemory_714 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  DMemory_715 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  DMemory_716 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  DMemory_717 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  DMemory_718 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  DMemory_719 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  DMemory_720 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  DMemory_721 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  DMemory_722 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  DMemory_723 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  DMemory_724 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  DMemory_725 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  DMemory_726 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  DMemory_727 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  DMemory_728 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  DMemory_729 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  DMemory_730 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  DMemory_731 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  DMemory_732 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  DMemory_733 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  DMemory_734 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  DMemory_735 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  DMemory_736 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  DMemory_737 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  DMemory_738 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  DMemory_739 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  DMemory_740 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  DMemory_741 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  DMemory_742 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  DMemory_743 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  DMemory_744 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  DMemory_745 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  DMemory_746 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  DMemory_747 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  DMemory_748 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  DMemory_749 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  DMemory_750 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  DMemory_751 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  DMemory_752 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  DMemory_753 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  DMemory_754 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  DMemory_755 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  DMemory_756 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  DMemory_757 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  DMemory_758 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  DMemory_759 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  DMemory_760 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  DMemory_761 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  DMemory_762 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  DMemory_763 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  DMemory_764 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  DMemory_765 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  DMemory_766 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  DMemory_767 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  DMemory_768 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  DMemory_769 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  DMemory_770 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  DMemory_771 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  DMemory_772 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  DMemory_773 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  DMemory_774 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  DMemory_775 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  DMemory_776 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  DMemory_777 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  DMemory_778 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  DMemory_779 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  DMemory_780 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  DMemory_781 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  DMemory_782 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  DMemory_783 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  DMemory_784 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  DMemory_785 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  DMemory_786 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  DMemory_787 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  DMemory_788 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  DMemory_789 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  DMemory_790 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  DMemory_791 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  DMemory_792 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  DMemory_793 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  DMemory_794 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  DMemory_795 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  DMemory_796 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  DMemory_797 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  DMemory_798 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  DMemory_799 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  DMemory_800 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  DMemory_801 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  DMemory_802 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  DMemory_803 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  DMemory_804 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  DMemory_805 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  DMemory_806 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  DMemory_807 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  DMemory_808 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  DMemory_809 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  DMemory_810 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  DMemory_811 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  DMemory_812 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  DMemory_813 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  DMemory_814 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  DMemory_815 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  DMemory_816 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  DMemory_817 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  DMemory_818 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  DMemory_819 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  DMemory_820 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  DMemory_821 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  DMemory_822 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  DMemory_823 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  DMemory_824 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  DMemory_825 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  DMemory_826 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  DMemory_827 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  DMemory_828 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  DMemory_829 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  DMemory_830 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  DMemory_831 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  DMemory_832 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  DMemory_833 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  DMemory_834 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  DMemory_835 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  DMemory_836 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  DMemory_837 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  DMemory_838 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  DMemory_839 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  DMemory_840 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  DMemory_841 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  DMemory_842 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  DMemory_843 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  DMemory_844 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  DMemory_845 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  DMemory_846 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  DMemory_847 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  DMemory_848 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  DMemory_849 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  DMemory_850 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  DMemory_851 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  DMemory_852 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  DMemory_853 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  DMemory_854 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  DMemory_855 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  DMemory_856 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  DMemory_857 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  DMemory_858 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  DMemory_859 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  DMemory_860 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  DMemory_861 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  DMemory_862 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  DMemory_863 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  DMemory_864 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  DMemory_865 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  DMemory_866 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  DMemory_867 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  DMemory_868 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  DMemory_869 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  DMemory_870 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  DMemory_871 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  DMemory_872 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  DMemory_873 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  DMemory_874 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  DMemory_875 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  DMemory_876 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  DMemory_877 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  DMemory_878 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  DMemory_879 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  DMemory_880 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  DMemory_881 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  DMemory_882 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  DMemory_883 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  DMemory_884 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  DMemory_885 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  DMemory_886 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  DMemory_887 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  DMemory_888 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  DMemory_889 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  DMemory_890 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  DMemory_891 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  DMemory_892 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  DMemory_893 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  DMemory_894 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  DMemory_895 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  DMemory_896 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  DMemory_897 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  DMemory_898 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  DMemory_899 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  DMemory_900 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  DMemory_901 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  DMemory_902 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  DMemory_903 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  DMemory_904 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  DMemory_905 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  DMemory_906 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  DMemory_907 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  DMemory_908 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  DMemory_909 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  DMemory_910 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  DMemory_911 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  DMemory_912 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  DMemory_913 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  DMemory_914 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  DMemory_915 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  DMemory_916 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  DMemory_917 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  DMemory_918 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  DMemory_919 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  DMemory_920 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  DMemory_921 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  DMemory_922 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  DMemory_923 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  DMemory_924 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  DMemory_925 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  DMemory_926 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  DMemory_927 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  DMemory_928 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  DMemory_929 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  DMemory_930 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  DMemory_931 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  DMemory_932 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  DMemory_933 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  DMemory_934 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  DMemory_935 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  DMemory_936 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  DMemory_937 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  DMemory_938 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  DMemory_939 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  DMemory_940 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  DMemory_941 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  DMemory_942 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  DMemory_943 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  DMemory_944 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  DMemory_945 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  DMemory_946 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  DMemory_947 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  DMemory_948 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  DMemory_949 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  DMemory_950 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  DMemory_951 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  DMemory_952 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  DMemory_953 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  DMemory_954 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  DMemory_955 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  DMemory_956 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  DMemory_957 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  DMemory_958 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  DMemory_959 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  DMemory_960 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  DMemory_961 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  DMemory_962 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  DMemory_963 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  DMemory_964 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  DMemory_965 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  DMemory_966 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  DMemory_967 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  DMemory_968 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  DMemory_969 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  DMemory_970 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  DMemory_971 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  DMemory_972 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  DMemory_973 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  DMemory_974 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  DMemory_975 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  DMemory_976 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  DMemory_977 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  DMemory_978 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  DMemory_979 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  DMemory_980 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  DMemory_981 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  DMemory_982 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  DMemory_983 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  DMemory_984 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  DMemory_985 = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  DMemory_986 = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  DMemory_987 = _RAND_1025[31:0];
  _RAND_1026 = {1{`RANDOM}};
  DMemory_988 = _RAND_1026[31:0];
  _RAND_1027 = {1{`RANDOM}};
  DMemory_989 = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  DMemory_990 = _RAND_1028[31:0];
  _RAND_1029 = {1{`RANDOM}};
  DMemory_991 = _RAND_1029[31:0];
  _RAND_1030 = {1{`RANDOM}};
  DMemory_992 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  DMemory_993 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  DMemory_994 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  DMemory_995 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  DMemory_996 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  DMemory_997 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  DMemory_998 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  DMemory_999 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  DMemory_1000 = _RAND_1038[31:0];
  _RAND_1039 = {1{`RANDOM}};
  DMemory_1001 = _RAND_1039[31:0];
  _RAND_1040 = {1{`RANDOM}};
  DMemory_1002 = _RAND_1040[31:0];
  _RAND_1041 = {1{`RANDOM}};
  DMemory_1003 = _RAND_1041[31:0];
  _RAND_1042 = {1{`RANDOM}};
  DMemory_1004 = _RAND_1042[31:0];
  _RAND_1043 = {1{`RANDOM}};
  DMemory_1005 = _RAND_1043[31:0];
  _RAND_1044 = {1{`RANDOM}};
  DMemory_1006 = _RAND_1044[31:0];
  _RAND_1045 = {1{`RANDOM}};
  DMemory_1007 = _RAND_1045[31:0];
  _RAND_1046 = {1{`RANDOM}};
  DMemory_1008 = _RAND_1046[31:0];
  _RAND_1047 = {1{`RANDOM}};
  DMemory_1009 = _RAND_1047[31:0];
  _RAND_1048 = {1{`RANDOM}};
  DMemory_1010 = _RAND_1048[31:0];
  _RAND_1049 = {1{`RANDOM}};
  DMemory_1011 = _RAND_1049[31:0];
  _RAND_1050 = {1{`RANDOM}};
  DMemory_1012 = _RAND_1050[31:0];
  _RAND_1051 = {1{`RANDOM}};
  DMemory_1013 = _RAND_1051[31:0];
  _RAND_1052 = {1{`RANDOM}};
  DMemory_1014 = _RAND_1052[31:0];
  _RAND_1053 = {1{`RANDOM}};
  DMemory_1015 = _RAND_1053[31:0];
  _RAND_1054 = {1{`RANDOM}};
  DMemory_1016 = _RAND_1054[31:0];
  _RAND_1055 = {1{`RANDOM}};
  DMemory_1017 = _RAND_1055[31:0];
  _RAND_1056 = {1{`RANDOM}};
  DMemory_1018 = _RAND_1056[31:0];
  _RAND_1057 = {1{`RANDOM}};
  DMemory_1019 = _RAND_1057[31:0];
  _RAND_1058 = {1{`RANDOM}};
  DMemory_1020 = _RAND_1058[31:0];
  _RAND_1059 = {1{`RANDOM}};
  DMemory_1021 = _RAND_1059[31:0];
  _RAND_1060 = {1{`RANDOM}};
  DMemory_1022 = _RAND_1060[31:0];
  _RAND_1061 = {1{`RANDOM}};
  DMemory_1023 = _RAND_1061[31:0];
  _RAND_1062 = {1{`RANDOM}};
  IMemory_0 = _RAND_1062[31:0];
  _RAND_1063 = {1{`RANDOM}};
  IMemory_1 = _RAND_1063[31:0];
  _RAND_1064 = {1{`RANDOM}};
  IMemory_2 = _RAND_1064[31:0];
  _RAND_1065 = {1{`RANDOM}};
  IMemory_3 = _RAND_1065[31:0];
  _RAND_1066 = {1{`RANDOM}};
  IFIDIR = _RAND_1066[31:0];
  _RAND_1067 = {1{`RANDOM}};
  IDEXIR = _RAND_1067[31:0];
  _RAND_1068 = {1{`RANDOM}};
  EXMEMIR = _RAND_1068[31:0];
  _RAND_1069 = {1{`RANDOM}};
  MEMWBIR = _RAND_1069[31:0];
  _RAND_1070 = {2{`RANDOM}};
  CurPC = _RAND_1070[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
