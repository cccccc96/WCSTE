module CAMCell(
  input   clock,
  input   reset,
  input   io_write,
  input   io_ki,
  input   io_di,
  output  io_lhi
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  oi; // @[cam.scala 15:19]
  wire  ti = io_write & io_di | ~io_write & oi; // @[cam.scala 17:29]
  assign io_lhi = oi & io_ki | ~oi & ~io_ki; // @[cam.scala 20:27]
  always @(posedge clock) begin
    if (reset) begin // @[cam.scala 15:19]
      oi <= 1'h0; // @[cam.scala 15:19]
    end else begin
      oi <= ti; // @[cam.scala 18:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  oi = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CAMLine_m(
  input         clock,
  input         reset,
  input         io_we,
  input         io_wi,
  input  [63:0] io_key,
  input  [63:0] io_din,
  output        io_hit
);
  wire  CAMCell_clock; // @[cam.scala 114:44]
  wire  CAMCell_reset; // @[cam.scala 114:44]
  wire  CAMCell_io_write; // @[cam.scala 114:44]
  wire  CAMCell_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_io_di; // @[cam.scala 114:44]
  wire  CAMCell_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_1_clock; // @[cam.scala 114:44]
  wire  CAMCell_1_reset; // @[cam.scala 114:44]
  wire  CAMCell_1_io_write; // @[cam.scala 114:44]
  wire  CAMCell_1_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_1_io_di; // @[cam.scala 114:44]
  wire  CAMCell_1_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_2_clock; // @[cam.scala 114:44]
  wire  CAMCell_2_reset; // @[cam.scala 114:44]
  wire  CAMCell_2_io_write; // @[cam.scala 114:44]
  wire  CAMCell_2_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_2_io_di; // @[cam.scala 114:44]
  wire  CAMCell_2_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_3_clock; // @[cam.scala 114:44]
  wire  CAMCell_3_reset; // @[cam.scala 114:44]
  wire  CAMCell_3_io_write; // @[cam.scala 114:44]
  wire  CAMCell_3_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_3_io_di; // @[cam.scala 114:44]
  wire  CAMCell_3_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_4_clock; // @[cam.scala 114:44]
  wire  CAMCell_4_reset; // @[cam.scala 114:44]
  wire  CAMCell_4_io_write; // @[cam.scala 114:44]
  wire  CAMCell_4_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_4_io_di; // @[cam.scala 114:44]
  wire  CAMCell_4_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_5_clock; // @[cam.scala 114:44]
  wire  CAMCell_5_reset; // @[cam.scala 114:44]
  wire  CAMCell_5_io_write; // @[cam.scala 114:44]
  wire  CAMCell_5_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_5_io_di; // @[cam.scala 114:44]
  wire  CAMCell_5_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_6_clock; // @[cam.scala 114:44]
  wire  CAMCell_6_reset; // @[cam.scala 114:44]
  wire  CAMCell_6_io_write; // @[cam.scala 114:44]
  wire  CAMCell_6_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_6_io_di; // @[cam.scala 114:44]
  wire  CAMCell_6_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_7_clock; // @[cam.scala 114:44]
  wire  CAMCell_7_reset; // @[cam.scala 114:44]
  wire  CAMCell_7_io_write; // @[cam.scala 114:44]
  wire  CAMCell_7_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_7_io_di; // @[cam.scala 114:44]
  wire  CAMCell_7_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_8_clock; // @[cam.scala 114:44]
  wire  CAMCell_8_reset; // @[cam.scala 114:44]
  wire  CAMCell_8_io_write; // @[cam.scala 114:44]
  wire  CAMCell_8_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_8_io_di; // @[cam.scala 114:44]
  wire  CAMCell_8_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_9_clock; // @[cam.scala 114:44]
  wire  CAMCell_9_reset; // @[cam.scala 114:44]
  wire  CAMCell_9_io_write; // @[cam.scala 114:44]
  wire  CAMCell_9_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_9_io_di; // @[cam.scala 114:44]
  wire  CAMCell_9_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_10_clock; // @[cam.scala 114:44]
  wire  CAMCell_10_reset; // @[cam.scala 114:44]
  wire  CAMCell_10_io_write; // @[cam.scala 114:44]
  wire  CAMCell_10_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_10_io_di; // @[cam.scala 114:44]
  wire  CAMCell_10_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_11_clock; // @[cam.scala 114:44]
  wire  CAMCell_11_reset; // @[cam.scala 114:44]
  wire  CAMCell_11_io_write; // @[cam.scala 114:44]
  wire  CAMCell_11_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_11_io_di; // @[cam.scala 114:44]
  wire  CAMCell_11_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_12_clock; // @[cam.scala 114:44]
  wire  CAMCell_12_reset; // @[cam.scala 114:44]
  wire  CAMCell_12_io_write; // @[cam.scala 114:44]
  wire  CAMCell_12_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_12_io_di; // @[cam.scala 114:44]
  wire  CAMCell_12_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_13_clock; // @[cam.scala 114:44]
  wire  CAMCell_13_reset; // @[cam.scala 114:44]
  wire  CAMCell_13_io_write; // @[cam.scala 114:44]
  wire  CAMCell_13_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_13_io_di; // @[cam.scala 114:44]
  wire  CAMCell_13_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_14_clock; // @[cam.scala 114:44]
  wire  CAMCell_14_reset; // @[cam.scala 114:44]
  wire  CAMCell_14_io_write; // @[cam.scala 114:44]
  wire  CAMCell_14_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_14_io_di; // @[cam.scala 114:44]
  wire  CAMCell_14_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_15_clock; // @[cam.scala 114:44]
  wire  CAMCell_15_reset; // @[cam.scala 114:44]
  wire  CAMCell_15_io_write; // @[cam.scala 114:44]
  wire  CAMCell_15_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_15_io_di; // @[cam.scala 114:44]
  wire  CAMCell_15_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_16_clock; // @[cam.scala 114:44]
  wire  CAMCell_16_reset; // @[cam.scala 114:44]
  wire  CAMCell_16_io_write; // @[cam.scala 114:44]
  wire  CAMCell_16_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_16_io_di; // @[cam.scala 114:44]
  wire  CAMCell_16_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_17_clock; // @[cam.scala 114:44]
  wire  CAMCell_17_reset; // @[cam.scala 114:44]
  wire  CAMCell_17_io_write; // @[cam.scala 114:44]
  wire  CAMCell_17_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_17_io_di; // @[cam.scala 114:44]
  wire  CAMCell_17_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_18_clock; // @[cam.scala 114:44]
  wire  CAMCell_18_reset; // @[cam.scala 114:44]
  wire  CAMCell_18_io_write; // @[cam.scala 114:44]
  wire  CAMCell_18_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_18_io_di; // @[cam.scala 114:44]
  wire  CAMCell_18_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_19_clock; // @[cam.scala 114:44]
  wire  CAMCell_19_reset; // @[cam.scala 114:44]
  wire  CAMCell_19_io_write; // @[cam.scala 114:44]
  wire  CAMCell_19_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_19_io_di; // @[cam.scala 114:44]
  wire  CAMCell_19_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_20_clock; // @[cam.scala 114:44]
  wire  CAMCell_20_reset; // @[cam.scala 114:44]
  wire  CAMCell_20_io_write; // @[cam.scala 114:44]
  wire  CAMCell_20_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_20_io_di; // @[cam.scala 114:44]
  wire  CAMCell_20_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_21_clock; // @[cam.scala 114:44]
  wire  CAMCell_21_reset; // @[cam.scala 114:44]
  wire  CAMCell_21_io_write; // @[cam.scala 114:44]
  wire  CAMCell_21_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_21_io_di; // @[cam.scala 114:44]
  wire  CAMCell_21_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_22_clock; // @[cam.scala 114:44]
  wire  CAMCell_22_reset; // @[cam.scala 114:44]
  wire  CAMCell_22_io_write; // @[cam.scala 114:44]
  wire  CAMCell_22_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_22_io_di; // @[cam.scala 114:44]
  wire  CAMCell_22_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_23_clock; // @[cam.scala 114:44]
  wire  CAMCell_23_reset; // @[cam.scala 114:44]
  wire  CAMCell_23_io_write; // @[cam.scala 114:44]
  wire  CAMCell_23_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_23_io_di; // @[cam.scala 114:44]
  wire  CAMCell_23_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_24_clock; // @[cam.scala 114:44]
  wire  CAMCell_24_reset; // @[cam.scala 114:44]
  wire  CAMCell_24_io_write; // @[cam.scala 114:44]
  wire  CAMCell_24_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_24_io_di; // @[cam.scala 114:44]
  wire  CAMCell_24_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_25_clock; // @[cam.scala 114:44]
  wire  CAMCell_25_reset; // @[cam.scala 114:44]
  wire  CAMCell_25_io_write; // @[cam.scala 114:44]
  wire  CAMCell_25_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_25_io_di; // @[cam.scala 114:44]
  wire  CAMCell_25_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_26_clock; // @[cam.scala 114:44]
  wire  CAMCell_26_reset; // @[cam.scala 114:44]
  wire  CAMCell_26_io_write; // @[cam.scala 114:44]
  wire  CAMCell_26_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_26_io_di; // @[cam.scala 114:44]
  wire  CAMCell_26_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_27_clock; // @[cam.scala 114:44]
  wire  CAMCell_27_reset; // @[cam.scala 114:44]
  wire  CAMCell_27_io_write; // @[cam.scala 114:44]
  wire  CAMCell_27_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_27_io_di; // @[cam.scala 114:44]
  wire  CAMCell_27_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_28_clock; // @[cam.scala 114:44]
  wire  CAMCell_28_reset; // @[cam.scala 114:44]
  wire  CAMCell_28_io_write; // @[cam.scala 114:44]
  wire  CAMCell_28_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_28_io_di; // @[cam.scala 114:44]
  wire  CAMCell_28_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_29_clock; // @[cam.scala 114:44]
  wire  CAMCell_29_reset; // @[cam.scala 114:44]
  wire  CAMCell_29_io_write; // @[cam.scala 114:44]
  wire  CAMCell_29_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_29_io_di; // @[cam.scala 114:44]
  wire  CAMCell_29_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_30_clock; // @[cam.scala 114:44]
  wire  CAMCell_30_reset; // @[cam.scala 114:44]
  wire  CAMCell_30_io_write; // @[cam.scala 114:44]
  wire  CAMCell_30_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_30_io_di; // @[cam.scala 114:44]
  wire  CAMCell_30_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_31_clock; // @[cam.scala 114:44]
  wire  CAMCell_31_reset; // @[cam.scala 114:44]
  wire  CAMCell_31_io_write; // @[cam.scala 114:44]
  wire  CAMCell_31_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_31_io_di; // @[cam.scala 114:44]
  wire  CAMCell_31_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_32_clock; // @[cam.scala 114:44]
  wire  CAMCell_32_reset; // @[cam.scala 114:44]
  wire  CAMCell_32_io_write; // @[cam.scala 114:44]
  wire  CAMCell_32_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_32_io_di; // @[cam.scala 114:44]
  wire  CAMCell_32_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_33_clock; // @[cam.scala 114:44]
  wire  CAMCell_33_reset; // @[cam.scala 114:44]
  wire  CAMCell_33_io_write; // @[cam.scala 114:44]
  wire  CAMCell_33_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_33_io_di; // @[cam.scala 114:44]
  wire  CAMCell_33_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_34_clock; // @[cam.scala 114:44]
  wire  CAMCell_34_reset; // @[cam.scala 114:44]
  wire  CAMCell_34_io_write; // @[cam.scala 114:44]
  wire  CAMCell_34_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_34_io_di; // @[cam.scala 114:44]
  wire  CAMCell_34_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_35_clock; // @[cam.scala 114:44]
  wire  CAMCell_35_reset; // @[cam.scala 114:44]
  wire  CAMCell_35_io_write; // @[cam.scala 114:44]
  wire  CAMCell_35_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_35_io_di; // @[cam.scala 114:44]
  wire  CAMCell_35_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_36_clock; // @[cam.scala 114:44]
  wire  CAMCell_36_reset; // @[cam.scala 114:44]
  wire  CAMCell_36_io_write; // @[cam.scala 114:44]
  wire  CAMCell_36_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_36_io_di; // @[cam.scala 114:44]
  wire  CAMCell_36_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_37_clock; // @[cam.scala 114:44]
  wire  CAMCell_37_reset; // @[cam.scala 114:44]
  wire  CAMCell_37_io_write; // @[cam.scala 114:44]
  wire  CAMCell_37_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_37_io_di; // @[cam.scala 114:44]
  wire  CAMCell_37_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_38_clock; // @[cam.scala 114:44]
  wire  CAMCell_38_reset; // @[cam.scala 114:44]
  wire  CAMCell_38_io_write; // @[cam.scala 114:44]
  wire  CAMCell_38_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_38_io_di; // @[cam.scala 114:44]
  wire  CAMCell_38_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_39_clock; // @[cam.scala 114:44]
  wire  CAMCell_39_reset; // @[cam.scala 114:44]
  wire  CAMCell_39_io_write; // @[cam.scala 114:44]
  wire  CAMCell_39_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_39_io_di; // @[cam.scala 114:44]
  wire  CAMCell_39_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_40_clock; // @[cam.scala 114:44]
  wire  CAMCell_40_reset; // @[cam.scala 114:44]
  wire  CAMCell_40_io_write; // @[cam.scala 114:44]
  wire  CAMCell_40_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_40_io_di; // @[cam.scala 114:44]
  wire  CAMCell_40_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_41_clock; // @[cam.scala 114:44]
  wire  CAMCell_41_reset; // @[cam.scala 114:44]
  wire  CAMCell_41_io_write; // @[cam.scala 114:44]
  wire  CAMCell_41_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_41_io_di; // @[cam.scala 114:44]
  wire  CAMCell_41_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_42_clock; // @[cam.scala 114:44]
  wire  CAMCell_42_reset; // @[cam.scala 114:44]
  wire  CAMCell_42_io_write; // @[cam.scala 114:44]
  wire  CAMCell_42_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_42_io_di; // @[cam.scala 114:44]
  wire  CAMCell_42_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_43_clock; // @[cam.scala 114:44]
  wire  CAMCell_43_reset; // @[cam.scala 114:44]
  wire  CAMCell_43_io_write; // @[cam.scala 114:44]
  wire  CAMCell_43_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_43_io_di; // @[cam.scala 114:44]
  wire  CAMCell_43_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_44_clock; // @[cam.scala 114:44]
  wire  CAMCell_44_reset; // @[cam.scala 114:44]
  wire  CAMCell_44_io_write; // @[cam.scala 114:44]
  wire  CAMCell_44_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_44_io_di; // @[cam.scala 114:44]
  wire  CAMCell_44_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_45_clock; // @[cam.scala 114:44]
  wire  CAMCell_45_reset; // @[cam.scala 114:44]
  wire  CAMCell_45_io_write; // @[cam.scala 114:44]
  wire  CAMCell_45_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_45_io_di; // @[cam.scala 114:44]
  wire  CAMCell_45_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_46_clock; // @[cam.scala 114:44]
  wire  CAMCell_46_reset; // @[cam.scala 114:44]
  wire  CAMCell_46_io_write; // @[cam.scala 114:44]
  wire  CAMCell_46_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_46_io_di; // @[cam.scala 114:44]
  wire  CAMCell_46_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_47_clock; // @[cam.scala 114:44]
  wire  CAMCell_47_reset; // @[cam.scala 114:44]
  wire  CAMCell_47_io_write; // @[cam.scala 114:44]
  wire  CAMCell_47_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_47_io_di; // @[cam.scala 114:44]
  wire  CAMCell_47_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_48_clock; // @[cam.scala 114:44]
  wire  CAMCell_48_reset; // @[cam.scala 114:44]
  wire  CAMCell_48_io_write; // @[cam.scala 114:44]
  wire  CAMCell_48_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_48_io_di; // @[cam.scala 114:44]
  wire  CAMCell_48_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_49_clock; // @[cam.scala 114:44]
  wire  CAMCell_49_reset; // @[cam.scala 114:44]
  wire  CAMCell_49_io_write; // @[cam.scala 114:44]
  wire  CAMCell_49_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_49_io_di; // @[cam.scala 114:44]
  wire  CAMCell_49_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_50_clock; // @[cam.scala 114:44]
  wire  CAMCell_50_reset; // @[cam.scala 114:44]
  wire  CAMCell_50_io_write; // @[cam.scala 114:44]
  wire  CAMCell_50_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_50_io_di; // @[cam.scala 114:44]
  wire  CAMCell_50_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_51_clock; // @[cam.scala 114:44]
  wire  CAMCell_51_reset; // @[cam.scala 114:44]
  wire  CAMCell_51_io_write; // @[cam.scala 114:44]
  wire  CAMCell_51_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_51_io_di; // @[cam.scala 114:44]
  wire  CAMCell_51_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_52_clock; // @[cam.scala 114:44]
  wire  CAMCell_52_reset; // @[cam.scala 114:44]
  wire  CAMCell_52_io_write; // @[cam.scala 114:44]
  wire  CAMCell_52_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_52_io_di; // @[cam.scala 114:44]
  wire  CAMCell_52_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_53_clock; // @[cam.scala 114:44]
  wire  CAMCell_53_reset; // @[cam.scala 114:44]
  wire  CAMCell_53_io_write; // @[cam.scala 114:44]
  wire  CAMCell_53_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_53_io_di; // @[cam.scala 114:44]
  wire  CAMCell_53_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_54_clock; // @[cam.scala 114:44]
  wire  CAMCell_54_reset; // @[cam.scala 114:44]
  wire  CAMCell_54_io_write; // @[cam.scala 114:44]
  wire  CAMCell_54_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_54_io_di; // @[cam.scala 114:44]
  wire  CAMCell_54_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_55_clock; // @[cam.scala 114:44]
  wire  CAMCell_55_reset; // @[cam.scala 114:44]
  wire  CAMCell_55_io_write; // @[cam.scala 114:44]
  wire  CAMCell_55_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_55_io_di; // @[cam.scala 114:44]
  wire  CAMCell_55_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_56_clock; // @[cam.scala 114:44]
  wire  CAMCell_56_reset; // @[cam.scala 114:44]
  wire  CAMCell_56_io_write; // @[cam.scala 114:44]
  wire  CAMCell_56_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_56_io_di; // @[cam.scala 114:44]
  wire  CAMCell_56_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_57_clock; // @[cam.scala 114:44]
  wire  CAMCell_57_reset; // @[cam.scala 114:44]
  wire  CAMCell_57_io_write; // @[cam.scala 114:44]
  wire  CAMCell_57_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_57_io_di; // @[cam.scala 114:44]
  wire  CAMCell_57_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_58_clock; // @[cam.scala 114:44]
  wire  CAMCell_58_reset; // @[cam.scala 114:44]
  wire  CAMCell_58_io_write; // @[cam.scala 114:44]
  wire  CAMCell_58_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_58_io_di; // @[cam.scala 114:44]
  wire  CAMCell_58_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_59_clock; // @[cam.scala 114:44]
  wire  CAMCell_59_reset; // @[cam.scala 114:44]
  wire  CAMCell_59_io_write; // @[cam.scala 114:44]
  wire  CAMCell_59_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_59_io_di; // @[cam.scala 114:44]
  wire  CAMCell_59_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_60_clock; // @[cam.scala 114:44]
  wire  CAMCell_60_reset; // @[cam.scala 114:44]
  wire  CAMCell_60_io_write; // @[cam.scala 114:44]
  wire  CAMCell_60_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_60_io_di; // @[cam.scala 114:44]
  wire  CAMCell_60_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_61_clock; // @[cam.scala 114:44]
  wire  CAMCell_61_reset; // @[cam.scala 114:44]
  wire  CAMCell_61_io_write; // @[cam.scala 114:44]
  wire  CAMCell_61_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_61_io_di; // @[cam.scala 114:44]
  wire  CAMCell_61_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_62_clock; // @[cam.scala 114:44]
  wire  CAMCell_62_reset; // @[cam.scala 114:44]
  wire  CAMCell_62_io_write; // @[cam.scala 114:44]
  wire  CAMCell_62_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_62_io_di; // @[cam.scala 114:44]
  wire  CAMCell_62_io_lhi; // @[cam.scala 114:44]
  wire  CAMCell_63_clock; // @[cam.scala 114:44]
  wire  CAMCell_63_reset; // @[cam.scala 114:44]
  wire  CAMCell_63_io_write; // @[cam.scala 114:44]
  wire  CAMCell_63_io_ki; // @[cam.scala 114:44]
  wire  CAMCell_63_io_di; // @[cam.scala 114:44]
  wire  CAMCell_63_io_lhi; // @[cam.scala 114:44]
  wire  camCells_0_lhi = CAMCell_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_1_lhi = CAMCell_1_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_2_lhi = CAMCell_2_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_3_lhi = CAMCell_3_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_4_lhi = CAMCell_4_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_5_lhi = CAMCell_5_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_6_lhi = CAMCell_6_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_7_lhi = CAMCell_7_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_8_lhi = CAMCell_8_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_9_lhi = CAMCell_9_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_10_lhi = CAMCell_10_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_11_lhi = CAMCell_11_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_12_lhi = CAMCell_12_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_13_lhi = CAMCell_13_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_14_lhi = CAMCell_14_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_15_lhi = CAMCell_15_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_16_lhi = CAMCell_16_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_17_lhi = CAMCell_17_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_18_lhi = CAMCell_18_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_19_lhi = CAMCell_19_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_20_lhi = CAMCell_20_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_21_lhi = CAMCell_21_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_22_lhi = CAMCell_22_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_23_lhi = CAMCell_23_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_24_lhi = CAMCell_24_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_25_lhi = CAMCell_25_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_26_lhi = CAMCell_26_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_27_lhi = CAMCell_27_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_28_lhi = CAMCell_28_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_29_lhi = CAMCell_29_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_30_lhi = CAMCell_30_io_lhi; // @[cam.scala 114:{25,25}]
  wire  _io_hit_T_29 = camCells_0_lhi & camCells_1_lhi & camCells_2_lhi & camCells_3_lhi & camCells_4_lhi &
    camCells_5_lhi & camCells_6_lhi & camCells_7_lhi & camCells_8_lhi & camCells_9_lhi & camCells_10_lhi &
    camCells_11_lhi & camCells_12_lhi & camCells_13_lhi & camCells_14_lhi & camCells_15_lhi & camCells_16_lhi &
    camCells_17_lhi & camCells_18_lhi & camCells_19_lhi & camCells_20_lhi & camCells_21_lhi & camCells_22_lhi &
    camCells_23_lhi & camCells_24_lhi & camCells_25_lhi & camCells_26_lhi & camCells_27_lhi & camCells_28_lhi &
    camCells_29_lhi & camCells_30_lhi; // @[cam.scala 123:27]
  wire  camCells_31_lhi = CAMCell_31_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_32_lhi = CAMCell_32_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_33_lhi = CAMCell_33_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_34_lhi = CAMCell_34_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_35_lhi = CAMCell_35_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_36_lhi = CAMCell_36_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_37_lhi = CAMCell_37_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_38_lhi = CAMCell_38_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_39_lhi = CAMCell_39_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_40_lhi = CAMCell_40_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_41_lhi = CAMCell_41_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_42_lhi = CAMCell_42_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_43_lhi = CAMCell_43_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_44_lhi = CAMCell_44_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_45_lhi = CAMCell_45_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_46_lhi = CAMCell_46_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_47_lhi = CAMCell_47_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_48_lhi = CAMCell_48_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_49_lhi = CAMCell_49_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_50_lhi = CAMCell_50_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_51_lhi = CAMCell_51_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_52_lhi = CAMCell_52_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_53_lhi = CAMCell_53_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_54_lhi = CAMCell_54_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_55_lhi = CAMCell_55_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_56_lhi = CAMCell_56_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_57_lhi = CAMCell_57_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_58_lhi = CAMCell_58_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_59_lhi = CAMCell_59_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_60_lhi = CAMCell_60_io_lhi; // @[cam.scala 114:{25,25}]
  wire  _io_hit_T_59 = _io_hit_T_29 & camCells_31_lhi & camCells_32_lhi & camCells_33_lhi & camCells_34_lhi &
    camCells_35_lhi & camCells_36_lhi & camCells_37_lhi & camCells_38_lhi & camCells_39_lhi & camCells_40_lhi &
    camCells_41_lhi & camCells_42_lhi & camCells_43_lhi & camCells_44_lhi & camCells_45_lhi & camCells_46_lhi &
    camCells_47_lhi & camCells_48_lhi & camCells_49_lhi & camCells_50_lhi & camCells_51_lhi & camCells_52_lhi &
    camCells_53_lhi & camCells_54_lhi & camCells_55_lhi & camCells_56_lhi & camCells_57_lhi & camCells_58_lhi &
    camCells_59_lhi & camCells_60_lhi; // @[cam.scala 123:27]
  wire  camCells_61_lhi = CAMCell_61_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_62_lhi = CAMCell_62_io_lhi; // @[cam.scala 114:{25,25}]
  wire  camCells_63_lhi = CAMCell_63_io_lhi; // @[cam.scala 114:{25,25}]
  CAMCell CAMCell ( // @[cam.scala 114:44]
    .clock(CAMCell_clock),
    .reset(CAMCell_reset),
    .io_write(CAMCell_io_write),
    .io_ki(CAMCell_io_ki),
    .io_di(CAMCell_io_di),
    .io_lhi(CAMCell_io_lhi)
  );
  CAMCell CAMCell_1 ( // @[cam.scala 114:44]
    .clock(CAMCell_1_clock),
    .reset(CAMCell_1_reset),
    .io_write(CAMCell_1_io_write),
    .io_ki(CAMCell_1_io_ki),
    .io_di(CAMCell_1_io_di),
    .io_lhi(CAMCell_1_io_lhi)
  );
  CAMCell CAMCell_2 ( // @[cam.scala 114:44]
    .clock(CAMCell_2_clock),
    .reset(CAMCell_2_reset),
    .io_write(CAMCell_2_io_write),
    .io_ki(CAMCell_2_io_ki),
    .io_di(CAMCell_2_io_di),
    .io_lhi(CAMCell_2_io_lhi)
  );
  CAMCell CAMCell_3 ( // @[cam.scala 114:44]
    .clock(CAMCell_3_clock),
    .reset(CAMCell_3_reset),
    .io_write(CAMCell_3_io_write),
    .io_ki(CAMCell_3_io_ki),
    .io_di(CAMCell_3_io_di),
    .io_lhi(CAMCell_3_io_lhi)
  );
  CAMCell CAMCell_4 ( // @[cam.scala 114:44]
    .clock(CAMCell_4_clock),
    .reset(CAMCell_4_reset),
    .io_write(CAMCell_4_io_write),
    .io_ki(CAMCell_4_io_ki),
    .io_di(CAMCell_4_io_di),
    .io_lhi(CAMCell_4_io_lhi)
  );
  CAMCell CAMCell_5 ( // @[cam.scala 114:44]
    .clock(CAMCell_5_clock),
    .reset(CAMCell_5_reset),
    .io_write(CAMCell_5_io_write),
    .io_ki(CAMCell_5_io_ki),
    .io_di(CAMCell_5_io_di),
    .io_lhi(CAMCell_5_io_lhi)
  );
  CAMCell CAMCell_6 ( // @[cam.scala 114:44]
    .clock(CAMCell_6_clock),
    .reset(CAMCell_6_reset),
    .io_write(CAMCell_6_io_write),
    .io_ki(CAMCell_6_io_ki),
    .io_di(CAMCell_6_io_di),
    .io_lhi(CAMCell_6_io_lhi)
  );
  CAMCell CAMCell_7 ( // @[cam.scala 114:44]
    .clock(CAMCell_7_clock),
    .reset(CAMCell_7_reset),
    .io_write(CAMCell_7_io_write),
    .io_ki(CAMCell_7_io_ki),
    .io_di(CAMCell_7_io_di),
    .io_lhi(CAMCell_7_io_lhi)
  );
  CAMCell CAMCell_8 ( // @[cam.scala 114:44]
    .clock(CAMCell_8_clock),
    .reset(CAMCell_8_reset),
    .io_write(CAMCell_8_io_write),
    .io_ki(CAMCell_8_io_ki),
    .io_di(CAMCell_8_io_di),
    .io_lhi(CAMCell_8_io_lhi)
  );
  CAMCell CAMCell_9 ( // @[cam.scala 114:44]
    .clock(CAMCell_9_clock),
    .reset(CAMCell_9_reset),
    .io_write(CAMCell_9_io_write),
    .io_ki(CAMCell_9_io_ki),
    .io_di(CAMCell_9_io_di),
    .io_lhi(CAMCell_9_io_lhi)
  );
  CAMCell CAMCell_10 ( // @[cam.scala 114:44]
    .clock(CAMCell_10_clock),
    .reset(CAMCell_10_reset),
    .io_write(CAMCell_10_io_write),
    .io_ki(CAMCell_10_io_ki),
    .io_di(CAMCell_10_io_di),
    .io_lhi(CAMCell_10_io_lhi)
  );
  CAMCell CAMCell_11 ( // @[cam.scala 114:44]
    .clock(CAMCell_11_clock),
    .reset(CAMCell_11_reset),
    .io_write(CAMCell_11_io_write),
    .io_ki(CAMCell_11_io_ki),
    .io_di(CAMCell_11_io_di),
    .io_lhi(CAMCell_11_io_lhi)
  );
  CAMCell CAMCell_12 ( // @[cam.scala 114:44]
    .clock(CAMCell_12_clock),
    .reset(CAMCell_12_reset),
    .io_write(CAMCell_12_io_write),
    .io_ki(CAMCell_12_io_ki),
    .io_di(CAMCell_12_io_di),
    .io_lhi(CAMCell_12_io_lhi)
  );
  CAMCell CAMCell_13 ( // @[cam.scala 114:44]
    .clock(CAMCell_13_clock),
    .reset(CAMCell_13_reset),
    .io_write(CAMCell_13_io_write),
    .io_ki(CAMCell_13_io_ki),
    .io_di(CAMCell_13_io_di),
    .io_lhi(CAMCell_13_io_lhi)
  );
  CAMCell CAMCell_14 ( // @[cam.scala 114:44]
    .clock(CAMCell_14_clock),
    .reset(CAMCell_14_reset),
    .io_write(CAMCell_14_io_write),
    .io_ki(CAMCell_14_io_ki),
    .io_di(CAMCell_14_io_di),
    .io_lhi(CAMCell_14_io_lhi)
  );
  CAMCell CAMCell_15 ( // @[cam.scala 114:44]
    .clock(CAMCell_15_clock),
    .reset(CAMCell_15_reset),
    .io_write(CAMCell_15_io_write),
    .io_ki(CAMCell_15_io_ki),
    .io_di(CAMCell_15_io_di),
    .io_lhi(CAMCell_15_io_lhi)
  );
  CAMCell CAMCell_16 ( // @[cam.scala 114:44]
    .clock(CAMCell_16_clock),
    .reset(CAMCell_16_reset),
    .io_write(CAMCell_16_io_write),
    .io_ki(CAMCell_16_io_ki),
    .io_di(CAMCell_16_io_di),
    .io_lhi(CAMCell_16_io_lhi)
  );
  CAMCell CAMCell_17 ( // @[cam.scala 114:44]
    .clock(CAMCell_17_clock),
    .reset(CAMCell_17_reset),
    .io_write(CAMCell_17_io_write),
    .io_ki(CAMCell_17_io_ki),
    .io_di(CAMCell_17_io_di),
    .io_lhi(CAMCell_17_io_lhi)
  );
  CAMCell CAMCell_18 ( // @[cam.scala 114:44]
    .clock(CAMCell_18_clock),
    .reset(CAMCell_18_reset),
    .io_write(CAMCell_18_io_write),
    .io_ki(CAMCell_18_io_ki),
    .io_di(CAMCell_18_io_di),
    .io_lhi(CAMCell_18_io_lhi)
  );
  CAMCell CAMCell_19 ( // @[cam.scala 114:44]
    .clock(CAMCell_19_clock),
    .reset(CAMCell_19_reset),
    .io_write(CAMCell_19_io_write),
    .io_ki(CAMCell_19_io_ki),
    .io_di(CAMCell_19_io_di),
    .io_lhi(CAMCell_19_io_lhi)
  );
  CAMCell CAMCell_20 ( // @[cam.scala 114:44]
    .clock(CAMCell_20_clock),
    .reset(CAMCell_20_reset),
    .io_write(CAMCell_20_io_write),
    .io_ki(CAMCell_20_io_ki),
    .io_di(CAMCell_20_io_di),
    .io_lhi(CAMCell_20_io_lhi)
  );
  CAMCell CAMCell_21 ( // @[cam.scala 114:44]
    .clock(CAMCell_21_clock),
    .reset(CAMCell_21_reset),
    .io_write(CAMCell_21_io_write),
    .io_ki(CAMCell_21_io_ki),
    .io_di(CAMCell_21_io_di),
    .io_lhi(CAMCell_21_io_lhi)
  );
  CAMCell CAMCell_22 ( // @[cam.scala 114:44]
    .clock(CAMCell_22_clock),
    .reset(CAMCell_22_reset),
    .io_write(CAMCell_22_io_write),
    .io_ki(CAMCell_22_io_ki),
    .io_di(CAMCell_22_io_di),
    .io_lhi(CAMCell_22_io_lhi)
  );
  CAMCell CAMCell_23 ( // @[cam.scala 114:44]
    .clock(CAMCell_23_clock),
    .reset(CAMCell_23_reset),
    .io_write(CAMCell_23_io_write),
    .io_ki(CAMCell_23_io_ki),
    .io_di(CAMCell_23_io_di),
    .io_lhi(CAMCell_23_io_lhi)
  );
  CAMCell CAMCell_24 ( // @[cam.scala 114:44]
    .clock(CAMCell_24_clock),
    .reset(CAMCell_24_reset),
    .io_write(CAMCell_24_io_write),
    .io_ki(CAMCell_24_io_ki),
    .io_di(CAMCell_24_io_di),
    .io_lhi(CAMCell_24_io_lhi)
  );
  CAMCell CAMCell_25 ( // @[cam.scala 114:44]
    .clock(CAMCell_25_clock),
    .reset(CAMCell_25_reset),
    .io_write(CAMCell_25_io_write),
    .io_ki(CAMCell_25_io_ki),
    .io_di(CAMCell_25_io_di),
    .io_lhi(CAMCell_25_io_lhi)
  );
  CAMCell CAMCell_26 ( // @[cam.scala 114:44]
    .clock(CAMCell_26_clock),
    .reset(CAMCell_26_reset),
    .io_write(CAMCell_26_io_write),
    .io_ki(CAMCell_26_io_ki),
    .io_di(CAMCell_26_io_di),
    .io_lhi(CAMCell_26_io_lhi)
  );
  CAMCell CAMCell_27 ( // @[cam.scala 114:44]
    .clock(CAMCell_27_clock),
    .reset(CAMCell_27_reset),
    .io_write(CAMCell_27_io_write),
    .io_ki(CAMCell_27_io_ki),
    .io_di(CAMCell_27_io_di),
    .io_lhi(CAMCell_27_io_lhi)
  );
  CAMCell CAMCell_28 ( // @[cam.scala 114:44]
    .clock(CAMCell_28_clock),
    .reset(CAMCell_28_reset),
    .io_write(CAMCell_28_io_write),
    .io_ki(CAMCell_28_io_ki),
    .io_di(CAMCell_28_io_di),
    .io_lhi(CAMCell_28_io_lhi)
  );
  CAMCell CAMCell_29 ( // @[cam.scala 114:44]
    .clock(CAMCell_29_clock),
    .reset(CAMCell_29_reset),
    .io_write(CAMCell_29_io_write),
    .io_ki(CAMCell_29_io_ki),
    .io_di(CAMCell_29_io_di),
    .io_lhi(CAMCell_29_io_lhi)
  );
  CAMCell CAMCell_30 ( // @[cam.scala 114:44]
    .clock(CAMCell_30_clock),
    .reset(CAMCell_30_reset),
    .io_write(CAMCell_30_io_write),
    .io_ki(CAMCell_30_io_ki),
    .io_di(CAMCell_30_io_di),
    .io_lhi(CAMCell_30_io_lhi)
  );
  CAMCell CAMCell_31 ( // @[cam.scala 114:44]
    .clock(CAMCell_31_clock),
    .reset(CAMCell_31_reset),
    .io_write(CAMCell_31_io_write),
    .io_ki(CAMCell_31_io_ki),
    .io_di(CAMCell_31_io_di),
    .io_lhi(CAMCell_31_io_lhi)
  );
  CAMCell CAMCell_32 ( // @[cam.scala 114:44]
    .clock(CAMCell_32_clock),
    .reset(CAMCell_32_reset),
    .io_write(CAMCell_32_io_write),
    .io_ki(CAMCell_32_io_ki),
    .io_di(CAMCell_32_io_di),
    .io_lhi(CAMCell_32_io_lhi)
  );
  CAMCell CAMCell_33 ( // @[cam.scala 114:44]
    .clock(CAMCell_33_clock),
    .reset(CAMCell_33_reset),
    .io_write(CAMCell_33_io_write),
    .io_ki(CAMCell_33_io_ki),
    .io_di(CAMCell_33_io_di),
    .io_lhi(CAMCell_33_io_lhi)
  );
  CAMCell CAMCell_34 ( // @[cam.scala 114:44]
    .clock(CAMCell_34_clock),
    .reset(CAMCell_34_reset),
    .io_write(CAMCell_34_io_write),
    .io_ki(CAMCell_34_io_ki),
    .io_di(CAMCell_34_io_di),
    .io_lhi(CAMCell_34_io_lhi)
  );
  CAMCell CAMCell_35 ( // @[cam.scala 114:44]
    .clock(CAMCell_35_clock),
    .reset(CAMCell_35_reset),
    .io_write(CAMCell_35_io_write),
    .io_ki(CAMCell_35_io_ki),
    .io_di(CAMCell_35_io_di),
    .io_lhi(CAMCell_35_io_lhi)
  );
  CAMCell CAMCell_36 ( // @[cam.scala 114:44]
    .clock(CAMCell_36_clock),
    .reset(CAMCell_36_reset),
    .io_write(CAMCell_36_io_write),
    .io_ki(CAMCell_36_io_ki),
    .io_di(CAMCell_36_io_di),
    .io_lhi(CAMCell_36_io_lhi)
  );
  CAMCell CAMCell_37 ( // @[cam.scala 114:44]
    .clock(CAMCell_37_clock),
    .reset(CAMCell_37_reset),
    .io_write(CAMCell_37_io_write),
    .io_ki(CAMCell_37_io_ki),
    .io_di(CAMCell_37_io_di),
    .io_lhi(CAMCell_37_io_lhi)
  );
  CAMCell CAMCell_38 ( // @[cam.scala 114:44]
    .clock(CAMCell_38_clock),
    .reset(CAMCell_38_reset),
    .io_write(CAMCell_38_io_write),
    .io_ki(CAMCell_38_io_ki),
    .io_di(CAMCell_38_io_di),
    .io_lhi(CAMCell_38_io_lhi)
  );
  CAMCell CAMCell_39 ( // @[cam.scala 114:44]
    .clock(CAMCell_39_clock),
    .reset(CAMCell_39_reset),
    .io_write(CAMCell_39_io_write),
    .io_ki(CAMCell_39_io_ki),
    .io_di(CAMCell_39_io_di),
    .io_lhi(CAMCell_39_io_lhi)
  );
  CAMCell CAMCell_40 ( // @[cam.scala 114:44]
    .clock(CAMCell_40_clock),
    .reset(CAMCell_40_reset),
    .io_write(CAMCell_40_io_write),
    .io_ki(CAMCell_40_io_ki),
    .io_di(CAMCell_40_io_di),
    .io_lhi(CAMCell_40_io_lhi)
  );
  CAMCell CAMCell_41 ( // @[cam.scala 114:44]
    .clock(CAMCell_41_clock),
    .reset(CAMCell_41_reset),
    .io_write(CAMCell_41_io_write),
    .io_ki(CAMCell_41_io_ki),
    .io_di(CAMCell_41_io_di),
    .io_lhi(CAMCell_41_io_lhi)
  );
  CAMCell CAMCell_42 ( // @[cam.scala 114:44]
    .clock(CAMCell_42_clock),
    .reset(CAMCell_42_reset),
    .io_write(CAMCell_42_io_write),
    .io_ki(CAMCell_42_io_ki),
    .io_di(CAMCell_42_io_di),
    .io_lhi(CAMCell_42_io_lhi)
  );
  CAMCell CAMCell_43 ( // @[cam.scala 114:44]
    .clock(CAMCell_43_clock),
    .reset(CAMCell_43_reset),
    .io_write(CAMCell_43_io_write),
    .io_ki(CAMCell_43_io_ki),
    .io_di(CAMCell_43_io_di),
    .io_lhi(CAMCell_43_io_lhi)
  );
  CAMCell CAMCell_44 ( // @[cam.scala 114:44]
    .clock(CAMCell_44_clock),
    .reset(CAMCell_44_reset),
    .io_write(CAMCell_44_io_write),
    .io_ki(CAMCell_44_io_ki),
    .io_di(CAMCell_44_io_di),
    .io_lhi(CAMCell_44_io_lhi)
  );
  CAMCell CAMCell_45 ( // @[cam.scala 114:44]
    .clock(CAMCell_45_clock),
    .reset(CAMCell_45_reset),
    .io_write(CAMCell_45_io_write),
    .io_ki(CAMCell_45_io_ki),
    .io_di(CAMCell_45_io_di),
    .io_lhi(CAMCell_45_io_lhi)
  );
  CAMCell CAMCell_46 ( // @[cam.scala 114:44]
    .clock(CAMCell_46_clock),
    .reset(CAMCell_46_reset),
    .io_write(CAMCell_46_io_write),
    .io_ki(CAMCell_46_io_ki),
    .io_di(CAMCell_46_io_di),
    .io_lhi(CAMCell_46_io_lhi)
  );
  CAMCell CAMCell_47 ( // @[cam.scala 114:44]
    .clock(CAMCell_47_clock),
    .reset(CAMCell_47_reset),
    .io_write(CAMCell_47_io_write),
    .io_ki(CAMCell_47_io_ki),
    .io_di(CAMCell_47_io_di),
    .io_lhi(CAMCell_47_io_lhi)
  );
  CAMCell CAMCell_48 ( // @[cam.scala 114:44]
    .clock(CAMCell_48_clock),
    .reset(CAMCell_48_reset),
    .io_write(CAMCell_48_io_write),
    .io_ki(CAMCell_48_io_ki),
    .io_di(CAMCell_48_io_di),
    .io_lhi(CAMCell_48_io_lhi)
  );
  CAMCell CAMCell_49 ( // @[cam.scala 114:44]
    .clock(CAMCell_49_clock),
    .reset(CAMCell_49_reset),
    .io_write(CAMCell_49_io_write),
    .io_ki(CAMCell_49_io_ki),
    .io_di(CAMCell_49_io_di),
    .io_lhi(CAMCell_49_io_lhi)
  );
  CAMCell CAMCell_50 ( // @[cam.scala 114:44]
    .clock(CAMCell_50_clock),
    .reset(CAMCell_50_reset),
    .io_write(CAMCell_50_io_write),
    .io_ki(CAMCell_50_io_ki),
    .io_di(CAMCell_50_io_di),
    .io_lhi(CAMCell_50_io_lhi)
  );
  CAMCell CAMCell_51 ( // @[cam.scala 114:44]
    .clock(CAMCell_51_clock),
    .reset(CAMCell_51_reset),
    .io_write(CAMCell_51_io_write),
    .io_ki(CAMCell_51_io_ki),
    .io_di(CAMCell_51_io_di),
    .io_lhi(CAMCell_51_io_lhi)
  );
  CAMCell CAMCell_52 ( // @[cam.scala 114:44]
    .clock(CAMCell_52_clock),
    .reset(CAMCell_52_reset),
    .io_write(CAMCell_52_io_write),
    .io_ki(CAMCell_52_io_ki),
    .io_di(CAMCell_52_io_di),
    .io_lhi(CAMCell_52_io_lhi)
  );
  CAMCell CAMCell_53 ( // @[cam.scala 114:44]
    .clock(CAMCell_53_clock),
    .reset(CAMCell_53_reset),
    .io_write(CAMCell_53_io_write),
    .io_ki(CAMCell_53_io_ki),
    .io_di(CAMCell_53_io_di),
    .io_lhi(CAMCell_53_io_lhi)
  );
  CAMCell CAMCell_54 ( // @[cam.scala 114:44]
    .clock(CAMCell_54_clock),
    .reset(CAMCell_54_reset),
    .io_write(CAMCell_54_io_write),
    .io_ki(CAMCell_54_io_ki),
    .io_di(CAMCell_54_io_di),
    .io_lhi(CAMCell_54_io_lhi)
  );
  CAMCell CAMCell_55 ( // @[cam.scala 114:44]
    .clock(CAMCell_55_clock),
    .reset(CAMCell_55_reset),
    .io_write(CAMCell_55_io_write),
    .io_ki(CAMCell_55_io_ki),
    .io_di(CAMCell_55_io_di),
    .io_lhi(CAMCell_55_io_lhi)
  );
  CAMCell CAMCell_56 ( // @[cam.scala 114:44]
    .clock(CAMCell_56_clock),
    .reset(CAMCell_56_reset),
    .io_write(CAMCell_56_io_write),
    .io_ki(CAMCell_56_io_ki),
    .io_di(CAMCell_56_io_di),
    .io_lhi(CAMCell_56_io_lhi)
  );
  CAMCell CAMCell_57 ( // @[cam.scala 114:44]
    .clock(CAMCell_57_clock),
    .reset(CAMCell_57_reset),
    .io_write(CAMCell_57_io_write),
    .io_ki(CAMCell_57_io_ki),
    .io_di(CAMCell_57_io_di),
    .io_lhi(CAMCell_57_io_lhi)
  );
  CAMCell CAMCell_58 ( // @[cam.scala 114:44]
    .clock(CAMCell_58_clock),
    .reset(CAMCell_58_reset),
    .io_write(CAMCell_58_io_write),
    .io_ki(CAMCell_58_io_ki),
    .io_di(CAMCell_58_io_di),
    .io_lhi(CAMCell_58_io_lhi)
  );
  CAMCell CAMCell_59 ( // @[cam.scala 114:44]
    .clock(CAMCell_59_clock),
    .reset(CAMCell_59_reset),
    .io_write(CAMCell_59_io_write),
    .io_ki(CAMCell_59_io_ki),
    .io_di(CAMCell_59_io_di),
    .io_lhi(CAMCell_59_io_lhi)
  );
  CAMCell CAMCell_60 ( // @[cam.scala 114:44]
    .clock(CAMCell_60_clock),
    .reset(CAMCell_60_reset),
    .io_write(CAMCell_60_io_write),
    .io_ki(CAMCell_60_io_ki),
    .io_di(CAMCell_60_io_di),
    .io_lhi(CAMCell_60_io_lhi)
  );
  CAMCell CAMCell_61 ( // @[cam.scala 114:44]
    .clock(CAMCell_61_clock),
    .reset(CAMCell_61_reset),
    .io_write(CAMCell_61_io_write),
    .io_ki(CAMCell_61_io_ki),
    .io_di(CAMCell_61_io_di),
    .io_lhi(CAMCell_61_io_lhi)
  );
  CAMCell CAMCell_62 ( // @[cam.scala 114:44]
    .clock(CAMCell_62_clock),
    .reset(CAMCell_62_reset),
    .io_write(CAMCell_62_io_write),
    .io_ki(CAMCell_62_io_ki),
    .io_di(CAMCell_62_io_di),
    .io_lhi(CAMCell_62_io_lhi)
  );
  CAMCell CAMCell_63 ( // @[cam.scala 114:44]
    .clock(CAMCell_63_clock),
    .reset(CAMCell_63_reset),
    .io_write(CAMCell_63_io_write),
    .io_ki(CAMCell_63_io_ki),
    .io_di(CAMCell_63_io_di),
    .io_lhi(CAMCell_63_io_lhi)
  );
  assign io_hit = _io_hit_T_59 & camCells_61_lhi & camCells_62_lhi & camCells_63_lhi; // @[cam.scala 123:27]
  assign CAMCell_clock = clock;
  assign CAMCell_reset = reset;
  assign CAMCell_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_io_ki = io_key[0]; // @[cam.scala 118:29]
  assign CAMCell_io_di = io_din[0]; // @[cam.scala 119:29]
  assign CAMCell_1_clock = clock;
  assign CAMCell_1_reset = reset;
  assign CAMCell_1_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_1_io_ki = io_key[1]; // @[cam.scala 118:29]
  assign CAMCell_1_io_di = io_din[1]; // @[cam.scala 119:29]
  assign CAMCell_2_clock = clock;
  assign CAMCell_2_reset = reset;
  assign CAMCell_2_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_2_io_ki = io_key[2]; // @[cam.scala 118:29]
  assign CAMCell_2_io_di = io_din[2]; // @[cam.scala 119:29]
  assign CAMCell_3_clock = clock;
  assign CAMCell_3_reset = reset;
  assign CAMCell_3_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_3_io_ki = io_key[3]; // @[cam.scala 118:29]
  assign CAMCell_3_io_di = io_din[3]; // @[cam.scala 119:29]
  assign CAMCell_4_clock = clock;
  assign CAMCell_4_reset = reset;
  assign CAMCell_4_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_4_io_ki = io_key[4]; // @[cam.scala 118:29]
  assign CAMCell_4_io_di = io_din[4]; // @[cam.scala 119:29]
  assign CAMCell_5_clock = clock;
  assign CAMCell_5_reset = reset;
  assign CAMCell_5_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_5_io_ki = io_key[5]; // @[cam.scala 118:29]
  assign CAMCell_5_io_di = io_din[5]; // @[cam.scala 119:29]
  assign CAMCell_6_clock = clock;
  assign CAMCell_6_reset = reset;
  assign CAMCell_6_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_6_io_ki = io_key[6]; // @[cam.scala 118:29]
  assign CAMCell_6_io_di = io_din[6]; // @[cam.scala 119:29]
  assign CAMCell_7_clock = clock;
  assign CAMCell_7_reset = reset;
  assign CAMCell_7_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_7_io_ki = io_key[7]; // @[cam.scala 118:29]
  assign CAMCell_7_io_di = io_din[7]; // @[cam.scala 119:29]
  assign CAMCell_8_clock = clock;
  assign CAMCell_8_reset = reset;
  assign CAMCell_8_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_8_io_ki = io_key[8]; // @[cam.scala 118:29]
  assign CAMCell_8_io_di = io_din[8]; // @[cam.scala 119:29]
  assign CAMCell_9_clock = clock;
  assign CAMCell_9_reset = reset;
  assign CAMCell_9_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_9_io_ki = io_key[9]; // @[cam.scala 118:29]
  assign CAMCell_9_io_di = io_din[9]; // @[cam.scala 119:29]
  assign CAMCell_10_clock = clock;
  assign CAMCell_10_reset = reset;
  assign CAMCell_10_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_10_io_ki = io_key[10]; // @[cam.scala 118:29]
  assign CAMCell_10_io_di = io_din[10]; // @[cam.scala 119:29]
  assign CAMCell_11_clock = clock;
  assign CAMCell_11_reset = reset;
  assign CAMCell_11_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_11_io_ki = io_key[11]; // @[cam.scala 118:29]
  assign CAMCell_11_io_di = io_din[11]; // @[cam.scala 119:29]
  assign CAMCell_12_clock = clock;
  assign CAMCell_12_reset = reset;
  assign CAMCell_12_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_12_io_ki = io_key[12]; // @[cam.scala 118:29]
  assign CAMCell_12_io_di = io_din[12]; // @[cam.scala 119:29]
  assign CAMCell_13_clock = clock;
  assign CAMCell_13_reset = reset;
  assign CAMCell_13_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_13_io_ki = io_key[13]; // @[cam.scala 118:29]
  assign CAMCell_13_io_di = io_din[13]; // @[cam.scala 119:29]
  assign CAMCell_14_clock = clock;
  assign CAMCell_14_reset = reset;
  assign CAMCell_14_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_14_io_ki = io_key[14]; // @[cam.scala 118:29]
  assign CAMCell_14_io_di = io_din[14]; // @[cam.scala 119:29]
  assign CAMCell_15_clock = clock;
  assign CAMCell_15_reset = reset;
  assign CAMCell_15_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_15_io_ki = io_key[15]; // @[cam.scala 118:29]
  assign CAMCell_15_io_di = io_din[15]; // @[cam.scala 119:29]
  assign CAMCell_16_clock = clock;
  assign CAMCell_16_reset = reset;
  assign CAMCell_16_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_16_io_ki = io_key[16]; // @[cam.scala 118:29]
  assign CAMCell_16_io_di = io_din[16]; // @[cam.scala 119:29]
  assign CAMCell_17_clock = clock;
  assign CAMCell_17_reset = reset;
  assign CAMCell_17_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_17_io_ki = io_key[17]; // @[cam.scala 118:29]
  assign CAMCell_17_io_di = io_din[17]; // @[cam.scala 119:29]
  assign CAMCell_18_clock = clock;
  assign CAMCell_18_reset = reset;
  assign CAMCell_18_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_18_io_ki = io_key[18]; // @[cam.scala 118:29]
  assign CAMCell_18_io_di = io_din[18]; // @[cam.scala 119:29]
  assign CAMCell_19_clock = clock;
  assign CAMCell_19_reset = reset;
  assign CAMCell_19_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_19_io_ki = io_key[19]; // @[cam.scala 118:29]
  assign CAMCell_19_io_di = io_din[19]; // @[cam.scala 119:29]
  assign CAMCell_20_clock = clock;
  assign CAMCell_20_reset = reset;
  assign CAMCell_20_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_20_io_ki = io_key[20]; // @[cam.scala 118:29]
  assign CAMCell_20_io_di = io_din[20]; // @[cam.scala 119:29]
  assign CAMCell_21_clock = clock;
  assign CAMCell_21_reset = reset;
  assign CAMCell_21_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_21_io_ki = io_key[21]; // @[cam.scala 118:29]
  assign CAMCell_21_io_di = io_din[21]; // @[cam.scala 119:29]
  assign CAMCell_22_clock = clock;
  assign CAMCell_22_reset = reset;
  assign CAMCell_22_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_22_io_ki = io_key[22]; // @[cam.scala 118:29]
  assign CAMCell_22_io_di = io_din[22]; // @[cam.scala 119:29]
  assign CAMCell_23_clock = clock;
  assign CAMCell_23_reset = reset;
  assign CAMCell_23_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_23_io_ki = io_key[23]; // @[cam.scala 118:29]
  assign CAMCell_23_io_di = io_din[23]; // @[cam.scala 119:29]
  assign CAMCell_24_clock = clock;
  assign CAMCell_24_reset = reset;
  assign CAMCell_24_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_24_io_ki = io_key[24]; // @[cam.scala 118:29]
  assign CAMCell_24_io_di = io_din[24]; // @[cam.scala 119:29]
  assign CAMCell_25_clock = clock;
  assign CAMCell_25_reset = reset;
  assign CAMCell_25_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_25_io_ki = io_key[25]; // @[cam.scala 118:29]
  assign CAMCell_25_io_di = io_din[25]; // @[cam.scala 119:29]
  assign CAMCell_26_clock = clock;
  assign CAMCell_26_reset = reset;
  assign CAMCell_26_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_26_io_ki = io_key[26]; // @[cam.scala 118:29]
  assign CAMCell_26_io_di = io_din[26]; // @[cam.scala 119:29]
  assign CAMCell_27_clock = clock;
  assign CAMCell_27_reset = reset;
  assign CAMCell_27_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_27_io_ki = io_key[27]; // @[cam.scala 118:29]
  assign CAMCell_27_io_di = io_din[27]; // @[cam.scala 119:29]
  assign CAMCell_28_clock = clock;
  assign CAMCell_28_reset = reset;
  assign CAMCell_28_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_28_io_ki = io_key[28]; // @[cam.scala 118:29]
  assign CAMCell_28_io_di = io_din[28]; // @[cam.scala 119:29]
  assign CAMCell_29_clock = clock;
  assign CAMCell_29_reset = reset;
  assign CAMCell_29_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_29_io_ki = io_key[29]; // @[cam.scala 118:29]
  assign CAMCell_29_io_di = io_din[29]; // @[cam.scala 119:29]
  assign CAMCell_30_clock = clock;
  assign CAMCell_30_reset = reset;
  assign CAMCell_30_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_30_io_ki = io_key[30]; // @[cam.scala 118:29]
  assign CAMCell_30_io_di = io_din[30]; // @[cam.scala 119:29]
  assign CAMCell_31_clock = clock;
  assign CAMCell_31_reset = reset;
  assign CAMCell_31_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_31_io_ki = io_key[31]; // @[cam.scala 118:29]
  assign CAMCell_31_io_di = io_din[31]; // @[cam.scala 119:29]
  assign CAMCell_32_clock = clock;
  assign CAMCell_32_reset = reset;
  assign CAMCell_32_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_32_io_ki = io_key[32]; // @[cam.scala 118:29]
  assign CAMCell_32_io_di = io_din[32]; // @[cam.scala 119:29]
  assign CAMCell_33_clock = clock;
  assign CAMCell_33_reset = reset;
  assign CAMCell_33_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_33_io_ki = io_key[33]; // @[cam.scala 118:29]
  assign CAMCell_33_io_di = io_din[33]; // @[cam.scala 119:29]
  assign CAMCell_34_clock = clock;
  assign CAMCell_34_reset = reset;
  assign CAMCell_34_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_34_io_ki = io_key[34]; // @[cam.scala 118:29]
  assign CAMCell_34_io_di = io_din[34]; // @[cam.scala 119:29]
  assign CAMCell_35_clock = clock;
  assign CAMCell_35_reset = reset;
  assign CAMCell_35_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_35_io_ki = io_key[35]; // @[cam.scala 118:29]
  assign CAMCell_35_io_di = io_din[35]; // @[cam.scala 119:29]
  assign CAMCell_36_clock = clock;
  assign CAMCell_36_reset = reset;
  assign CAMCell_36_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_36_io_ki = io_key[36]; // @[cam.scala 118:29]
  assign CAMCell_36_io_di = io_din[36]; // @[cam.scala 119:29]
  assign CAMCell_37_clock = clock;
  assign CAMCell_37_reset = reset;
  assign CAMCell_37_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_37_io_ki = io_key[37]; // @[cam.scala 118:29]
  assign CAMCell_37_io_di = io_din[37]; // @[cam.scala 119:29]
  assign CAMCell_38_clock = clock;
  assign CAMCell_38_reset = reset;
  assign CAMCell_38_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_38_io_ki = io_key[38]; // @[cam.scala 118:29]
  assign CAMCell_38_io_di = io_din[38]; // @[cam.scala 119:29]
  assign CAMCell_39_clock = clock;
  assign CAMCell_39_reset = reset;
  assign CAMCell_39_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_39_io_ki = io_key[39]; // @[cam.scala 118:29]
  assign CAMCell_39_io_di = io_din[39]; // @[cam.scala 119:29]
  assign CAMCell_40_clock = clock;
  assign CAMCell_40_reset = reset;
  assign CAMCell_40_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_40_io_ki = io_key[40]; // @[cam.scala 118:29]
  assign CAMCell_40_io_di = io_din[40]; // @[cam.scala 119:29]
  assign CAMCell_41_clock = clock;
  assign CAMCell_41_reset = reset;
  assign CAMCell_41_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_41_io_ki = io_key[41]; // @[cam.scala 118:29]
  assign CAMCell_41_io_di = io_din[41]; // @[cam.scala 119:29]
  assign CAMCell_42_clock = clock;
  assign CAMCell_42_reset = reset;
  assign CAMCell_42_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_42_io_ki = io_key[42]; // @[cam.scala 118:29]
  assign CAMCell_42_io_di = io_din[42]; // @[cam.scala 119:29]
  assign CAMCell_43_clock = clock;
  assign CAMCell_43_reset = reset;
  assign CAMCell_43_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_43_io_ki = io_key[43]; // @[cam.scala 118:29]
  assign CAMCell_43_io_di = io_din[43]; // @[cam.scala 119:29]
  assign CAMCell_44_clock = clock;
  assign CAMCell_44_reset = reset;
  assign CAMCell_44_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_44_io_ki = io_key[44]; // @[cam.scala 118:29]
  assign CAMCell_44_io_di = io_din[44]; // @[cam.scala 119:29]
  assign CAMCell_45_clock = clock;
  assign CAMCell_45_reset = reset;
  assign CAMCell_45_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_45_io_ki = io_key[45]; // @[cam.scala 118:29]
  assign CAMCell_45_io_di = io_din[45]; // @[cam.scala 119:29]
  assign CAMCell_46_clock = clock;
  assign CAMCell_46_reset = reset;
  assign CAMCell_46_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_46_io_ki = io_key[46]; // @[cam.scala 118:29]
  assign CAMCell_46_io_di = io_din[46]; // @[cam.scala 119:29]
  assign CAMCell_47_clock = clock;
  assign CAMCell_47_reset = reset;
  assign CAMCell_47_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_47_io_ki = io_key[47]; // @[cam.scala 118:29]
  assign CAMCell_47_io_di = io_din[47]; // @[cam.scala 119:29]
  assign CAMCell_48_clock = clock;
  assign CAMCell_48_reset = reset;
  assign CAMCell_48_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_48_io_ki = io_key[48]; // @[cam.scala 118:29]
  assign CAMCell_48_io_di = io_din[48]; // @[cam.scala 119:29]
  assign CAMCell_49_clock = clock;
  assign CAMCell_49_reset = reset;
  assign CAMCell_49_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_49_io_ki = io_key[49]; // @[cam.scala 118:29]
  assign CAMCell_49_io_di = io_din[49]; // @[cam.scala 119:29]
  assign CAMCell_50_clock = clock;
  assign CAMCell_50_reset = reset;
  assign CAMCell_50_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_50_io_ki = io_key[50]; // @[cam.scala 118:29]
  assign CAMCell_50_io_di = io_din[50]; // @[cam.scala 119:29]
  assign CAMCell_51_clock = clock;
  assign CAMCell_51_reset = reset;
  assign CAMCell_51_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_51_io_ki = io_key[51]; // @[cam.scala 118:29]
  assign CAMCell_51_io_di = io_din[51]; // @[cam.scala 119:29]
  assign CAMCell_52_clock = clock;
  assign CAMCell_52_reset = reset;
  assign CAMCell_52_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_52_io_ki = io_key[52]; // @[cam.scala 118:29]
  assign CAMCell_52_io_di = io_din[52]; // @[cam.scala 119:29]
  assign CAMCell_53_clock = clock;
  assign CAMCell_53_reset = reset;
  assign CAMCell_53_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_53_io_ki = io_key[53]; // @[cam.scala 118:29]
  assign CAMCell_53_io_di = io_din[53]; // @[cam.scala 119:29]
  assign CAMCell_54_clock = clock;
  assign CAMCell_54_reset = reset;
  assign CAMCell_54_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_54_io_ki = io_key[54]; // @[cam.scala 118:29]
  assign CAMCell_54_io_di = io_din[54]; // @[cam.scala 119:29]
  assign CAMCell_55_clock = clock;
  assign CAMCell_55_reset = reset;
  assign CAMCell_55_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_55_io_ki = io_key[55]; // @[cam.scala 118:29]
  assign CAMCell_55_io_di = io_din[55]; // @[cam.scala 119:29]
  assign CAMCell_56_clock = clock;
  assign CAMCell_56_reset = reset;
  assign CAMCell_56_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_56_io_ki = io_key[56]; // @[cam.scala 118:29]
  assign CAMCell_56_io_di = io_din[56]; // @[cam.scala 119:29]
  assign CAMCell_57_clock = clock;
  assign CAMCell_57_reset = reset;
  assign CAMCell_57_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_57_io_ki = io_key[57]; // @[cam.scala 118:29]
  assign CAMCell_57_io_di = io_din[57]; // @[cam.scala 119:29]
  assign CAMCell_58_clock = clock;
  assign CAMCell_58_reset = reset;
  assign CAMCell_58_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_58_io_ki = io_key[58]; // @[cam.scala 118:29]
  assign CAMCell_58_io_di = io_din[58]; // @[cam.scala 119:29]
  assign CAMCell_59_clock = clock;
  assign CAMCell_59_reset = reset;
  assign CAMCell_59_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_59_io_ki = io_key[59]; // @[cam.scala 118:29]
  assign CAMCell_59_io_di = io_din[59]; // @[cam.scala 119:29]
  assign CAMCell_60_clock = clock;
  assign CAMCell_60_reset = reset;
  assign CAMCell_60_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_60_io_ki = io_key[60]; // @[cam.scala 118:29]
  assign CAMCell_60_io_di = io_din[60]; // @[cam.scala 119:29]
  assign CAMCell_61_clock = clock;
  assign CAMCell_61_reset = reset;
  assign CAMCell_61_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_61_io_ki = io_key[61]; // @[cam.scala 118:29]
  assign CAMCell_61_io_di = io_din[61]; // @[cam.scala 119:29]
  assign CAMCell_62_clock = clock;
  assign CAMCell_62_reset = reset;
  assign CAMCell_62_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_62_io_ki = io_key[62]; // @[cam.scala 118:29]
  assign CAMCell_62_io_di = io_din[62]; // @[cam.scala 119:29]
  assign CAMCell_63_clock = clock;
  assign CAMCell_63_reset = reset;
  assign CAMCell_63_io_write = io_we & io_wi; // @[cam.scala 121:18]
  assign CAMCell_63_io_ki = io_key[63]; // @[cam.scala 118:29]
  assign CAMCell_63_io_di = io_din[63]; // @[cam.scala 119:29]
endmodule
module CAM_m_n(
  input         clock,
  input         reset,
  input         io_we,
  input  [63:0] io_key,
  input  [63:0] io_din,
  input  [63:0] io_waddr,
  output        io_hit
);
  wire  CAMLine_m_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_1_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_1_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_1_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_1_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_1_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_1_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_1_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_2_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_2_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_2_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_2_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_2_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_2_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_2_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_3_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_3_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_3_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_3_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_3_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_3_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_3_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_4_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_4_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_4_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_4_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_4_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_4_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_4_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_5_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_5_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_5_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_5_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_5_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_5_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_5_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_6_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_6_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_6_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_6_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_6_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_6_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_6_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_7_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_7_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_7_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_7_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_7_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_7_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_7_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_8_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_8_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_8_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_8_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_8_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_8_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_8_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_9_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_9_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_9_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_9_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_9_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_9_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_9_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_10_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_10_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_10_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_10_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_10_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_10_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_10_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_11_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_11_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_11_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_11_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_11_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_11_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_11_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_12_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_12_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_12_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_12_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_12_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_12_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_12_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_13_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_13_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_13_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_13_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_13_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_13_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_13_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_14_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_14_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_14_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_14_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_14_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_14_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_14_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_15_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_15_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_15_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_15_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_15_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_15_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_15_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_16_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_16_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_16_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_16_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_16_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_16_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_16_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_17_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_17_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_17_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_17_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_17_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_17_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_17_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_18_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_18_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_18_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_18_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_18_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_18_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_18_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_19_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_19_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_19_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_19_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_19_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_19_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_19_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_20_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_20_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_20_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_20_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_20_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_20_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_20_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_21_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_21_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_21_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_21_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_21_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_21_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_21_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_22_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_22_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_22_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_22_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_22_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_22_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_22_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_23_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_23_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_23_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_23_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_23_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_23_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_23_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_24_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_24_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_24_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_24_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_24_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_24_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_24_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_25_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_25_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_25_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_25_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_25_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_25_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_25_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_26_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_26_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_26_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_26_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_26_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_26_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_26_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_27_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_27_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_27_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_27_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_27_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_27_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_27_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_28_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_28_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_28_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_28_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_28_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_28_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_28_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_29_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_29_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_29_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_29_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_29_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_29_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_29_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_30_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_30_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_30_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_30_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_30_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_30_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_30_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_31_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_31_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_31_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_31_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_31_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_31_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_31_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_32_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_32_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_32_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_32_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_32_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_32_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_32_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_33_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_33_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_33_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_33_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_33_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_33_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_33_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_34_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_34_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_34_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_34_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_34_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_34_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_34_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_35_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_35_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_35_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_35_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_35_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_35_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_35_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_36_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_36_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_36_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_36_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_36_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_36_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_36_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_37_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_37_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_37_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_37_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_37_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_37_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_37_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_38_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_38_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_38_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_38_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_38_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_38_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_38_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_39_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_39_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_39_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_39_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_39_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_39_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_39_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_40_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_40_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_40_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_40_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_40_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_40_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_40_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_41_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_41_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_41_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_41_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_41_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_41_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_41_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_42_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_42_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_42_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_42_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_42_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_42_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_42_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_43_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_43_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_43_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_43_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_43_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_43_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_43_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_44_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_44_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_44_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_44_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_44_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_44_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_44_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_45_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_45_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_45_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_45_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_45_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_45_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_45_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_46_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_46_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_46_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_46_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_46_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_46_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_46_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_47_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_47_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_47_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_47_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_47_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_47_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_47_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_48_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_48_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_48_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_48_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_48_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_48_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_48_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_49_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_49_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_49_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_49_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_49_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_49_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_49_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_50_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_50_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_50_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_50_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_50_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_50_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_50_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_51_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_51_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_51_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_51_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_51_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_51_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_51_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_52_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_52_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_52_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_52_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_52_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_52_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_52_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_53_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_53_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_53_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_53_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_53_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_53_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_53_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_54_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_54_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_54_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_54_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_54_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_54_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_54_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_55_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_55_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_55_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_55_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_55_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_55_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_55_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_56_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_56_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_56_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_56_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_56_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_56_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_56_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_57_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_57_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_57_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_57_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_57_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_57_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_57_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_58_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_58_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_58_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_58_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_58_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_58_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_58_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_59_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_59_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_59_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_59_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_59_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_59_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_59_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_60_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_60_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_60_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_60_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_60_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_60_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_60_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_61_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_61_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_61_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_61_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_61_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_61_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_61_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_62_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_62_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_62_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_62_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_62_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_62_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_62_io_hit; // @[cam.scala 139:36]
  wire  CAMLine_m_63_clock; // @[cam.scala 139:36]
  wire  CAMLine_m_63_reset; // @[cam.scala 139:36]
  wire  CAMLine_m_63_io_we; // @[cam.scala 139:36]
  wire  CAMLine_m_63_io_wi; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_63_io_key; // @[cam.scala 139:36]
  wire [63:0] CAMLine_m_63_io_din; // @[cam.scala 139:36]
  wire  CAMLine_m_63_io_hit; // @[cam.scala 139:36]
  wire  _io_hit_T_29 = CAMLine_m_io_hit | CAMLine_m_1_io_hit | CAMLine_m_2_io_hit | CAMLine_m_3_io_hit |
    CAMLine_m_4_io_hit | CAMLine_m_5_io_hit | CAMLine_m_6_io_hit | CAMLine_m_7_io_hit | CAMLine_m_8_io_hit |
    CAMLine_m_9_io_hit | CAMLine_m_10_io_hit | CAMLine_m_11_io_hit | CAMLine_m_12_io_hit | CAMLine_m_13_io_hit |
    CAMLine_m_14_io_hit | CAMLine_m_15_io_hit | CAMLine_m_16_io_hit | CAMLine_m_17_io_hit | CAMLine_m_18_io_hit |
    CAMLine_m_19_io_hit | CAMLine_m_20_io_hit | CAMLine_m_21_io_hit | CAMLine_m_22_io_hit | CAMLine_m_23_io_hit |
    CAMLine_m_24_io_hit | CAMLine_m_25_io_hit | CAMLine_m_26_io_hit | CAMLine_m_27_io_hit | CAMLine_m_28_io_hit |
    CAMLine_m_29_io_hit | CAMLine_m_30_io_hit; // @[cam.scala 152:27]
  wire  _io_hit_T_59 = _io_hit_T_29 | CAMLine_m_31_io_hit | CAMLine_m_32_io_hit | CAMLine_m_33_io_hit |
    CAMLine_m_34_io_hit | CAMLine_m_35_io_hit | CAMLine_m_36_io_hit | CAMLine_m_37_io_hit | CAMLine_m_38_io_hit |
    CAMLine_m_39_io_hit | CAMLine_m_40_io_hit | CAMLine_m_41_io_hit | CAMLine_m_42_io_hit | CAMLine_m_43_io_hit |
    CAMLine_m_44_io_hit | CAMLine_m_45_io_hit | CAMLine_m_46_io_hit | CAMLine_m_47_io_hit | CAMLine_m_48_io_hit |
    CAMLine_m_49_io_hit | CAMLine_m_50_io_hit | CAMLine_m_51_io_hit | CAMLine_m_52_io_hit | CAMLine_m_53_io_hit |
    CAMLine_m_54_io_hit | CAMLine_m_55_io_hit | CAMLine_m_56_io_hit | CAMLine_m_57_io_hit | CAMLine_m_58_io_hit |
    CAMLine_m_59_io_hit | CAMLine_m_60_io_hit; // @[cam.scala 152:27]
  CAMLine_m CAMLine_m ( // @[cam.scala 139:36]
    .clock(CAMLine_m_clock),
    .reset(CAMLine_m_reset),
    .io_we(CAMLine_m_io_we),
    .io_wi(CAMLine_m_io_wi),
    .io_key(CAMLine_m_io_key),
    .io_din(CAMLine_m_io_din),
    .io_hit(CAMLine_m_io_hit)
  );
  CAMLine_m CAMLine_m_1 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_1_clock),
    .reset(CAMLine_m_1_reset),
    .io_we(CAMLine_m_1_io_we),
    .io_wi(CAMLine_m_1_io_wi),
    .io_key(CAMLine_m_1_io_key),
    .io_din(CAMLine_m_1_io_din),
    .io_hit(CAMLine_m_1_io_hit)
  );
  CAMLine_m CAMLine_m_2 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_2_clock),
    .reset(CAMLine_m_2_reset),
    .io_we(CAMLine_m_2_io_we),
    .io_wi(CAMLine_m_2_io_wi),
    .io_key(CAMLine_m_2_io_key),
    .io_din(CAMLine_m_2_io_din),
    .io_hit(CAMLine_m_2_io_hit)
  );
  CAMLine_m CAMLine_m_3 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_3_clock),
    .reset(CAMLine_m_3_reset),
    .io_we(CAMLine_m_3_io_we),
    .io_wi(CAMLine_m_3_io_wi),
    .io_key(CAMLine_m_3_io_key),
    .io_din(CAMLine_m_3_io_din),
    .io_hit(CAMLine_m_3_io_hit)
  );
  CAMLine_m CAMLine_m_4 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_4_clock),
    .reset(CAMLine_m_4_reset),
    .io_we(CAMLine_m_4_io_we),
    .io_wi(CAMLine_m_4_io_wi),
    .io_key(CAMLine_m_4_io_key),
    .io_din(CAMLine_m_4_io_din),
    .io_hit(CAMLine_m_4_io_hit)
  );
  CAMLine_m CAMLine_m_5 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_5_clock),
    .reset(CAMLine_m_5_reset),
    .io_we(CAMLine_m_5_io_we),
    .io_wi(CAMLine_m_5_io_wi),
    .io_key(CAMLine_m_5_io_key),
    .io_din(CAMLine_m_5_io_din),
    .io_hit(CAMLine_m_5_io_hit)
  );
  CAMLine_m CAMLine_m_6 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_6_clock),
    .reset(CAMLine_m_6_reset),
    .io_we(CAMLine_m_6_io_we),
    .io_wi(CAMLine_m_6_io_wi),
    .io_key(CAMLine_m_6_io_key),
    .io_din(CAMLine_m_6_io_din),
    .io_hit(CAMLine_m_6_io_hit)
  );
  CAMLine_m CAMLine_m_7 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_7_clock),
    .reset(CAMLine_m_7_reset),
    .io_we(CAMLine_m_7_io_we),
    .io_wi(CAMLine_m_7_io_wi),
    .io_key(CAMLine_m_7_io_key),
    .io_din(CAMLine_m_7_io_din),
    .io_hit(CAMLine_m_7_io_hit)
  );
  CAMLine_m CAMLine_m_8 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_8_clock),
    .reset(CAMLine_m_8_reset),
    .io_we(CAMLine_m_8_io_we),
    .io_wi(CAMLine_m_8_io_wi),
    .io_key(CAMLine_m_8_io_key),
    .io_din(CAMLine_m_8_io_din),
    .io_hit(CAMLine_m_8_io_hit)
  );
  CAMLine_m CAMLine_m_9 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_9_clock),
    .reset(CAMLine_m_9_reset),
    .io_we(CAMLine_m_9_io_we),
    .io_wi(CAMLine_m_9_io_wi),
    .io_key(CAMLine_m_9_io_key),
    .io_din(CAMLine_m_9_io_din),
    .io_hit(CAMLine_m_9_io_hit)
  );
  CAMLine_m CAMLine_m_10 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_10_clock),
    .reset(CAMLine_m_10_reset),
    .io_we(CAMLine_m_10_io_we),
    .io_wi(CAMLine_m_10_io_wi),
    .io_key(CAMLine_m_10_io_key),
    .io_din(CAMLine_m_10_io_din),
    .io_hit(CAMLine_m_10_io_hit)
  );
  CAMLine_m CAMLine_m_11 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_11_clock),
    .reset(CAMLine_m_11_reset),
    .io_we(CAMLine_m_11_io_we),
    .io_wi(CAMLine_m_11_io_wi),
    .io_key(CAMLine_m_11_io_key),
    .io_din(CAMLine_m_11_io_din),
    .io_hit(CAMLine_m_11_io_hit)
  );
  CAMLine_m CAMLine_m_12 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_12_clock),
    .reset(CAMLine_m_12_reset),
    .io_we(CAMLine_m_12_io_we),
    .io_wi(CAMLine_m_12_io_wi),
    .io_key(CAMLine_m_12_io_key),
    .io_din(CAMLine_m_12_io_din),
    .io_hit(CAMLine_m_12_io_hit)
  );
  CAMLine_m CAMLine_m_13 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_13_clock),
    .reset(CAMLine_m_13_reset),
    .io_we(CAMLine_m_13_io_we),
    .io_wi(CAMLine_m_13_io_wi),
    .io_key(CAMLine_m_13_io_key),
    .io_din(CAMLine_m_13_io_din),
    .io_hit(CAMLine_m_13_io_hit)
  );
  CAMLine_m CAMLine_m_14 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_14_clock),
    .reset(CAMLine_m_14_reset),
    .io_we(CAMLine_m_14_io_we),
    .io_wi(CAMLine_m_14_io_wi),
    .io_key(CAMLine_m_14_io_key),
    .io_din(CAMLine_m_14_io_din),
    .io_hit(CAMLine_m_14_io_hit)
  );
  CAMLine_m CAMLine_m_15 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_15_clock),
    .reset(CAMLine_m_15_reset),
    .io_we(CAMLine_m_15_io_we),
    .io_wi(CAMLine_m_15_io_wi),
    .io_key(CAMLine_m_15_io_key),
    .io_din(CAMLine_m_15_io_din),
    .io_hit(CAMLine_m_15_io_hit)
  );
  CAMLine_m CAMLine_m_16 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_16_clock),
    .reset(CAMLine_m_16_reset),
    .io_we(CAMLine_m_16_io_we),
    .io_wi(CAMLine_m_16_io_wi),
    .io_key(CAMLine_m_16_io_key),
    .io_din(CAMLine_m_16_io_din),
    .io_hit(CAMLine_m_16_io_hit)
  );
  CAMLine_m CAMLine_m_17 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_17_clock),
    .reset(CAMLine_m_17_reset),
    .io_we(CAMLine_m_17_io_we),
    .io_wi(CAMLine_m_17_io_wi),
    .io_key(CAMLine_m_17_io_key),
    .io_din(CAMLine_m_17_io_din),
    .io_hit(CAMLine_m_17_io_hit)
  );
  CAMLine_m CAMLine_m_18 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_18_clock),
    .reset(CAMLine_m_18_reset),
    .io_we(CAMLine_m_18_io_we),
    .io_wi(CAMLine_m_18_io_wi),
    .io_key(CAMLine_m_18_io_key),
    .io_din(CAMLine_m_18_io_din),
    .io_hit(CAMLine_m_18_io_hit)
  );
  CAMLine_m CAMLine_m_19 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_19_clock),
    .reset(CAMLine_m_19_reset),
    .io_we(CAMLine_m_19_io_we),
    .io_wi(CAMLine_m_19_io_wi),
    .io_key(CAMLine_m_19_io_key),
    .io_din(CAMLine_m_19_io_din),
    .io_hit(CAMLine_m_19_io_hit)
  );
  CAMLine_m CAMLine_m_20 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_20_clock),
    .reset(CAMLine_m_20_reset),
    .io_we(CAMLine_m_20_io_we),
    .io_wi(CAMLine_m_20_io_wi),
    .io_key(CAMLine_m_20_io_key),
    .io_din(CAMLine_m_20_io_din),
    .io_hit(CAMLine_m_20_io_hit)
  );
  CAMLine_m CAMLine_m_21 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_21_clock),
    .reset(CAMLine_m_21_reset),
    .io_we(CAMLine_m_21_io_we),
    .io_wi(CAMLine_m_21_io_wi),
    .io_key(CAMLine_m_21_io_key),
    .io_din(CAMLine_m_21_io_din),
    .io_hit(CAMLine_m_21_io_hit)
  );
  CAMLine_m CAMLine_m_22 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_22_clock),
    .reset(CAMLine_m_22_reset),
    .io_we(CAMLine_m_22_io_we),
    .io_wi(CAMLine_m_22_io_wi),
    .io_key(CAMLine_m_22_io_key),
    .io_din(CAMLine_m_22_io_din),
    .io_hit(CAMLine_m_22_io_hit)
  );
  CAMLine_m CAMLine_m_23 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_23_clock),
    .reset(CAMLine_m_23_reset),
    .io_we(CAMLine_m_23_io_we),
    .io_wi(CAMLine_m_23_io_wi),
    .io_key(CAMLine_m_23_io_key),
    .io_din(CAMLine_m_23_io_din),
    .io_hit(CAMLine_m_23_io_hit)
  );
  CAMLine_m CAMLine_m_24 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_24_clock),
    .reset(CAMLine_m_24_reset),
    .io_we(CAMLine_m_24_io_we),
    .io_wi(CAMLine_m_24_io_wi),
    .io_key(CAMLine_m_24_io_key),
    .io_din(CAMLine_m_24_io_din),
    .io_hit(CAMLine_m_24_io_hit)
  );
  CAMLine_m CAMLine_m_25 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_25_clock),
    .reset(CAMLine_m_25_reset),
    .io_we(CAMLine_m_25_io_we),
    .io_wi(CAMLine_m_25_io_wi),
    .io_key(CAMLine_m_25_io_key),
    .io_din(CAMLine_m_25_io_din),
    .io_hit(CAMLine_m_25_io_hit)
  );
  CAMLine_m CAMLine_m_26 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_26_clock),
    .reset(CAMLine_m_26_reset),
    .io_we(CAMLine_m_26_io_we),
    .io_wi(CAMLine_m_26_io_wi),
    .io_key(CAMLine_m_26_io_key),
    .io_din(CAMLine_m_26_io_din),
    .io_hit(CAMLine_m_26_io_hit)
  );
  CAMLine_m CAMLine_m_27 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_27_clock),
    .reset(CAMLine_m_27_reset),
    .io_we(CAMLine_m_27_io_we),
    .io_wi(CAMLine_m_27_io_wi),
    .io_key(CAMLine_m_27_io_key),
    .io_din(CAMLine_m_27_io_din),
    .io_hit(CAMLine_m_27_io_hit)
  );
  CAMLine_m CAMLine_m_28 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_28_clock),
    .reset(CAMLine_m_28_reset),
    .io_we(CAMLine_m_28_io_we),
    .io_wi(CAMLine_m_28_io_wi),
    .io_key(CAMLine_m_28_io_key),
    .io_din(CAMLine_m_28_io_din),
    .io_hit(CAMLine_m_28_io_hit)
  );
  CAMLine_m CAMLine_m_29 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_29_clock),
    .reset(CAMLine_m_29_reset),
    .io_we(CAMLine_m_29_io_we),
    .io_wi(CAMLine_m_29_io_wi),
    .io_key(CAMLine_m_29_io_key),
    .io_din(CAMLine_m_29_io_din),
    .io_hit(CAMLine_m_29_io_hit)
  );
  CAMLine_m CAMLine_m_30 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_30_clock),
    .reset(CAMLine_m_30_reset),
    .io_we(CAMLine_m_30_io_we),
    .io_wi(CAMLine_m_30_io_wi),
    .io_key(CAMLine_m_30_io_key),
    .io_din(CAMLine_m_30_io_din),
    .io_hit(CAMLine_m_30_io_hit)
  );
  CAMLine_m CAMLine_m_31 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_31_clock),
    .reset(CAMLine_m_31_reset),
    .io_we(CAMLine_m_31_io_we),
    .io_wi(CAMLine_m_31_io_wi),
    .io_key(CAMLine_m_31_io_key),
    .io_din(CAMLine_m_31_io_din),
    .io_hit(CAMLine_m_31_io_hit)
  );
  CAMLine_m CAMLine_m_32 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_32_clock),
    .reset(CAMLine_m_32_reset),
    .io_we(CAMLine_m_32_io_we),
    .io_wi(CAMLine_m_32_io_wi),
    .io_key(CAMLine_m_32_io_key),
    .io_din(CAMLine_m_32_io_din),
    .io_hit(CAMLine_m_32_io_hit)
  );
  CAMLine_m CAMLine_m_33 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_33_clock),
    .reset(CAMLine_m_33_reset),
    .io_we(CAMLine_m_33_io_we),
    .io_wi(CAMLine_m_33_io_wi),
    .io_key(CAMLine_m_33_io_key),
    .io_din(CAMLine_m_33_io_din),
    .io_hit(CAMLine_m_33_io_hit)
  );
  CAMLine_m CAMLine_m_34 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_34_clock),
    .reset(CAMLine_m_34_reset),
    .io_we(CAMLine_m_34_io_we),
    .io_wi(CAMLine_m_34_io_wi),
    .io_key(CAMLine_m_34_io_key),
    .io_din(CAMLine_m_34_io_din),
    .io_hit(CAMLine_m_34_io_hit)
  );
  CAMLine_m CAMLine_m_35 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_35_clock),
    .reset(CAMLine_m_35_reset),
    .io_we(CAMLine_m_35_io_we),
    .io_wi(CAMLine_m_35_io_wi),
    .io_key(CAMLine_m_35_io_key),
    .io_din(CAMLine_m_35_io_din),
    .io_hit(CAMLine_m_35_io_hit)
  );
  CAMLine_m CAMLine_m_36 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_36_clock),
    .reset(CAMLine_m_36_reset),
    .io_we(CAMLine_m_36_io_we),
    .io_wi(CAMLine_m_36_io_wi),
    .io_key(CAMLine_m_36_io_key),
    .io_din(CAMLine_m_36_io_din),
    .io_hit(CAMLine_m_36_io_hit)
  );
  CAMLine_m CAMLine_m_37 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_37_clock),
    .reset(CAMLine_m_37_reset),
    .io_we(CAMLine_m_37_io_we),
    .io_wi(CAMLine_m_37_io_wi),
    .io_key(CAMLine_m_37_io_key),
    .io_din(CAMLine_m_37_io_din),
    .io_hit(CAMLine_m_37_io_hit)
  );
  CAMLine_m CAMLine_m_38 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_38_clock),
    .reset(CAMLine_m_38_reset),
    .io_we(CAMLine_m_38_io_we),
    .io_wi(CAMLine_m_38_io_wi),
    .io_key(CAMLine_m_38_io_key),
    .io_din(CAMLine_m_38_io_din),
    .io_hit(CAMLine_m_38_io_hit)
  );
  CAMLine_m CAMLine_m_39 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_39_clock),
    .reset(CAMLine_m_39_reset),
    .io_we(CAMLine_m_39_io_we),
    .io_wi(CAMLine_m_39_io_wi),
    .io_key(CAMLine_m_39_io_key),
    .io_din(CAMLine_m_39_io_din),
    .io_hit(CAMLine_m_39_io_hit)
  );
  CAMLine_m CAMLine_m_40 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_40_clock),
    .reset(CAMLine_m_40_reset),
    .io_we(CAMLine_m_40_io_we),
    .io_wi(CAMLine_m_40_io_wi),
    .io_key(CAMLine_m_40_io_key),
    .io_din(CAMLine_m_40_io_din),
    .io_hit(CAMLine_m_40_io_hit)
  );
  CAMLine_m CAMLine_m_41 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_41_clock),
    .reset(CAMLine_m_41_reset),
    .io_we(CAMLine_m_41_io_we),
    .io_wi(CAMLine_m_41_io_wi),
    .io_key(CAMLine_m_41_io_key),
    .io_din(CAMLine_m_41_io_din),
    .io_hit(CAMLine_m_41_io_hit)
  );
  CAMLine_m CAMLine_m_42 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_42_clock),
    .reset(CAMLine_m_42_reset),
    .io_we(CAMLine_m_42_io_we),
    .io_wi(CAMLine_m_42_io_wi),
    .io_key(CAMLine_m_42_io_key),
    .io_din(CAMLine_m_42_io_din),
    .io_hit(CAMLine_m_42_io_hit)
  );
  CAMLine_m CAMLine_m_43 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_43_clock),
    .reset(CAMLine_m_43_reset),
    .io_we(CAMLine_m_43_io_we),
    .io_wi(CAMLine_m_43_io_wi),
    .io_key(CAMLine_m_43_io_key),
    .io_din(CAMLine_m_43_io_din),
    .io_hit(CAMLine_m_43_io_hit)
  );
  CAMLine_m CAMLine_m_44 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_44_clock),
    .reset(CAMLine_m_44_reset),
    .io_we(CAMLine_m_44_io_we),
    .io_wi(CAMLine_m_44_io_wi),
    .io_key(CAMLine_m_44_io_key),
    .io_din(CAMLine_m_44_io_din),
    .io_hit(CAMLine_m_44_io_hit)
  );
  CAMLine_m CAMLine_m_45 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_45_clock),
    .reset(CAMLine_m_45_reset),
    .io_we(CAMLine_m_45_io_we),
    .io_wi(CAMLine_m_45_io_wi),
    .io_key(CAMLine_m_45_io_key),
    .io_din(CAMLine_m_45_io_din),
    .io_hit(CAMLine_m_45_io_hit)
  );
  CAMLine_m CAMLine_m_46 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_46_clock),
    .reset(CAMLine_m_46_reset),
    .io_we(CAMLine_m_46_io_we),
    .io_wi(CAMLine_m_46_io_wi),
    .io_key(CAMLine_m_46_io_key),
    .io_din(CAMLine_m_46_io_din),
    .io_hit(CAMLine_m_46_io_hit)
  );
  CAMLine_m CAMLine_m_47 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_47_clock),
    .reset(CAMLine_m_47_reset),
    .io_we(CAMLine_m_47_io_we),
    .io_wi(CAMLine_m_47_io_wi),
    .io_key(CAMLine_m_47_io_key),
    .io_din(CAMLine_m_47_io_din),
    .io_hit(CAMLine_m_47_io_hit)
  );
  CAMLine_m CAMLine_m_48 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_48_clock),
    .reset(CAMLine_m_48_reset),
    .io_we(CAMLine_m_48_io_we),
    .io_wi(CAMLine_m_48_io_wi),
    .io_key(CAMLine_m_48_io_key),
    .io_din(CAMLine_m_48_io_din),
    .io_hit(CAMLine_m_48_io_hit)
  );
  CAMLine_m CAMLine_m_49 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_49_clock),
    .reset(CAMLine_m_49_reset),
    .io_we(CAMLine_m_49_io_we),
    .io_wi(CAMLine_m_49_io_wi),
    .io_key(CAMLine_m_49_io_key),
    .io_din(CAMLine_m_49_io_din),
    .io_hit(CAMLine_m_49_io_hit)
  );
  CAMLine_m CAMLine_m_50 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_50_clock),
    .reset(CAMLine_m_50_reset),
    .io_we(CAMLine_m_50_io_we),
    .io_wi(CAMLine_m_50_io_wi),
    .io_key(CAMLine_m_50_io_key),
    .io_din(CAMLine_m_50_io_din),
    .io_hit(CAMLine_m_50_io_hit)
  );
  CAMLine_m CAMLine_m_51 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_51_clock),
    .reset(CAMLine_m_51_reset),
    .io_we(CAMLine_m_51_io_we),
    .io_wi(CAMLine_m_51_io_wi),
    .io_key(CAMLine_m_51_io_key),
    .io_din(CAMLine_m_51_io_din),
    .io_hit(CAMLine_m_51_io_hit)
  );
  CAMLine_m CAMLine_m_52 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_52_clock),
    .reset(CAMLine_m_52_reset),
    .io_we(CAMLine_m_52_io_we),
    .io_wi(CAMLine_m_52_io_wi),
    .io_key(CAMLine_m_52_io_key),
    .io_din(CAMLine_m_52_io_din),
    .io_hit(CAMLine_m_52_io_hit)
  );
  CAMLine_m CAMLine_m_53 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_53_clock),
    .reset(CAMLine_m_53_reset),
    .io_we(CAMLine_m_53_io_we),
    .io_wi(CAMLine_m_53_io_wi),
    .io_key(CAMLine_m_53_io_key),
    .io_din(CAMLine_m_53_io_din),
    .io_hit(CAMLine_m_53_io_hit)
  );
  CAMLine_m CAMLine_m_54 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_54_clock),
    .reset(CAMLine_m_54_reset),
    .io_we(CAMLine_m_54_io_we),
    .io_wi(CAMLine_m_54_io_wi),
    .io_key(CAMLine_m_54_io_key),
    .io_din(CAMLine_m_54_io_din),
    .io_hit(CAMLine_m_54_io_hit)
  );
  CAMLine_m CAMLine_m_55 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_55_clock),
    .reset(CAMLine_m_55_reset),
    .io_we(CAMLine_m_55_io_we),
    .io_wi(CAMLine_m_55_io_wi),
    .io_key(CAMLine_m_55_io_key),
    .io_din(CAMLine_m_55_io_din),
    .io_hit(CAMLine_m_55_io_hit)
  );
  CAMLine_m CAMLine_m_56 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_56_clock),
    .reset(CAMLine_m_56_reset),
    .io_we(CAMLine_m_56_io_we),
    .io_wi(CAMLine_m_56_io_wi),
    .io_key(CAMLine_m_56_io_key),
    .io_din(CAMLine_m_56_io_din),
    .io_hit(CAMLine_m_56_io_hit)
  );
  CAMLine_m CAMLine_m_57 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_57_clock),
    .reset(CAMLine_m_57_reset),
    .io_we(CAMLine_m_57_io_we),
    .io_wi(CAMLine_m_57_io_wi),
    .io_key(CAMLine_m_57_io_key),
    .io_din(CAMLine_m_57_io_din),
    .io_hit(CAMLine_m_57_io_hit)
  );
  CAMLine_m CAMLine_m_58 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_58_clock),
    .reset(CAMLine_m_58_reset),
    .io_we(CAMLine_m_58_io_we),
    .io_wi(CAMLine_m_58_io_wi),
    .io_key(CAMLine_m_58_io_key),
    .io_din(CAMLine_m_58_io_din),
    .io_hit(CAMLine_m_58_io_hit)
  );
  CAMLine_m CAMLine_m_59 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_59_clock),
    .reset(CAMLine_m_59_reset),
    .io_we(CAMLine_m_59_io_we),
    .io_wi(CAMLine_m_59_io_wi),
    .io_key(CAMLine_m_59_io_key),
    .io_din(CAMLine_m_59_io_din),
    .io_hit(CAMLine_m_59_io_hit)
  );
  CAMLine_m CAMLine_m_60 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_60_clock),
    .reset(CAMLine_m_60_reset),
    .io_we(CAMLine_m_60_io_we),
    .io_wi(CAMLine_m_60_io_wi),
    .io_key(CAMLine_m_60_io_key),
    .io_din(CAMLine_m_60_io_din),
    .io_hit(CAMLine_m_60_io_hit)
  );
  CAMLine_m CAMLine_m_61 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_61_clock),
    .reset(CAMLine_m_61_reset),
    .io_we(CAMLine_m_61_io_we),
    .io_wi(CAMLine_m_61_io_wi),
    .io_key(CAMLine_m_61_io_key),
    .io_din(CAMLine_m_61_io_din),
    .io_hit(CAMLine_m_61_io_hit)
  );
  CAMLine_m CAMLine_m_62 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_62_clock),
    .reset(CAMLine_m_62_reset),
    .io_we(CAMLine_m_62_io_we),
    .io_wi(CAMLine_m_62_io_wi),
    .io_key(CAMLine_m_62_io_key),
    .io_din(CAMLine_m_62_io_din),
    .io_hit(CAMLine_m_62_io_hit)
  );
  CAMLine_m CAMLine_m_63 ( // @[cam.scala 139:36]
    .clock(CAMLine_m_63_clock),
    .reset(CAMLine_m_63_reset),
    .io_we(CAMLine_m_63_io_we),
    .io_wi(CAMLine_m_63_io_wi),
    .io_key(CAMLine_m_63_io_key),
    .io_din(CAMLine_m_63_io_din),
    .io_hit(CAMLine_m_63_io_hit)
  );
  assign io_hit = _io_hit_T_59 | CAMLine_m_61_io_hit | CAMLine_m_62_io_hit | CAMLine_m_63_io_hit; // @[cam.scala 152:27]
  assign CAMLine_m_clock = clock;
  assign CAMLine_m_reset = reset;
  assign CAMLine_m_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_io_wi = io_waddr[0]; // @[cam.scala 144:31]
  assign CAMLine_m_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_1_clock = clock;
  assign CAMLine_m_1_reset = reset;
  assign CAMLine_m_1_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_1_io_wi = io_waddr[1]; // @[cam.scala 144:31]
  assign CAMLine_m_1_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_1_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_2_clock = clock;
  assign CAMLine_m_2_reset = reset;
  assign CAMLine_m_2_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_2_io_wi = io_waddr[2]; // @[cam.scala 144:31]
  assign CAMLine_m_2_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_2_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_3_clock = clock;
  assign CAMLine_m_3_reset = reset;
  assign CAMLine_m_3_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_3_io_wi = io_waddr[3]; // @[cam.scala 144:31]
  assign CAMLine_m_3_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_3_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_4_clock = clock;
  assign CAMLine_m_4_reset = reset;
  assign CAMLine_m_4_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_4_io_wi = io_waddr[4]; // @[cam.scala 144:31]
  assign CAMLine_m_4_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_4_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_5_clock = clock;
  assign CAMLine_m_5_reset = reset;
  assign CAMLine_m_5_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_5_io_wi = io_waddr[5]; // @[cam.scala 144:31]
  assign CAMLine_m_5_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_5_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_6_clock = clock;
  assign CAMLine_m_6_reset = reset;
  assign CAMLine_m_6_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_6_io_wi = io_waddr[6]; // @[cam.scala 144:31]
  assign CAMLine_m_6_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_6_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_7_clock = clock;
  assign CAMLine_m_7_reset = reset;
  assign CAMLine_m_7_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_7_io_wi = io_waddr[7]; // @[cam.scala 144:31]
  assign CAMLine_m_7_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_7_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_8_clock = clock;
  assign CAMLine_m_8_reset = reset;
  assign CAMLine_m_8_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_8_io_wi = io_waddr[8]; // @[cam.scala 144:31]
  assign CAMLine_m_8_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_8_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_9_clock = clock;
  assign CAMLine_m_9_reset = reset;
  assign CAMLine_m_9_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_9_io_wi = io_waddr[9]; // @[cam.scala 144:31]
  assign CAMLine_m_9_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_9_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_10_clock = clock;
  assign CAMLine_m_10_reset = reset;
  assign CAMLine_m_10_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_10_io_wi = io_waddr[10]; // @[cam.scala 144:31]
  assign CAMLine_m_10_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_10_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_11_clock = clock;
  assign CAMLine_m_11_reset = reset;
  assign CAMLine_m_11_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_11_io_wi = io_waddr[11]; // @[cam.scala 144:31]
  assign CAMLine_m_11_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_11_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_12_clock = clock;
  assign CAMLine_m_12_reset = reset;
  assign CAMLine_m_12_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_12_io_wi = io_waddr[12]; // @[cam.scala 144:31]
  assign CAMLine_m_12_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_12_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_13_clock = clock;
  assign CAMLine_m_13_reset = reset;
  assign CAMLine_m_13_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_13_io_wi = io_waddr[13]; // @[cam.scala 144:31]
  assign CAMLine_m_13_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_13_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_14_clock = clock;
  assign CAMLine_m_14_reset = reset;
  assign CAMLine_m_14_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_14_io_wi = io_waddr[14]; // @[cam.scala 144:31]
  assign CAMLine_m_14_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_14_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_15_clock = clock;
  assign CAMLine_m_15_reset = reset;
  assign CAMLine_m_15_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_15_io_wi = io_waddr[15]; // @[cam.scala 144:31]
  assign CAMLine_m_15_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_15_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_16_clock = clock;
  assign CAMLine_m_16_reset = reset;
  assign CAMLine_m_16_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_16_io_wi = io_waddr[16]; // @[cam.scala 144:31]
  assign CAMLine_m_16_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_16_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_17_clock = clock;
  assign CAMLine_m_17_reset = reset;
  assign CAMLine_m_17_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_17_io_wi = io_waddr[17]; // @[cam.scala 144:31]
  assign CAMLine_m_17_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_17_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_18_clock = clock;
  assign CAMLine_m_18_reset = reset;
  assign CAMLine_m_18_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_18_io_wi = io_waddr[18]; // @[cam.scala 144:31]
  assign CAMLine_m_18_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_18_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_19_clock = clock;
  assign CAMLine_m_19_reset = reset;
  assign CAMLine_m_19_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_19_io_wi = io_waddr[19]; // @[cam.scala 144:31]
  assign CAMLine_m_19_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_19_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_20_clock = clock;
  assign CAMLine_m_20_reset = reset;
  assign CAMLine_m_20_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_20_io_wi = io_waddr[20]; // @[cam.scala 144:31]
  assign CAMLine_m_20_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_20_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_21_clock = clock;
  assign CAMLine_m_21_reset = reset;
  assign CAMLine_m_21_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_21_io_wi = io_waddr[21]; // @[cam.scala 144:31]
  assign CAMLine_m_21_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_21_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_22_clock = clock;
  assign CAMLine_m_22_reset = reset;
  assign CAMLine_m_22_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_22_io_wi = io_waddr[22]; // @[cam.scala 144:31]
  assign CAMLine_m_22_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_22_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_23_clock = clock;
  assign CAMLine_m_23_reset = reset;
  assign CAMLine_m_23_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_23_io_wi = io_waddr[23]; // @[cam.scala 144:31]
  assign CAMLine_m_23_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_23_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_24_clock = clock;
  assign CAMLine_m_24_reset = reset;
  assign CAMLine_m_24_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_24_io_wi = io_waddr[24]; // @[cam.scala 144:31]
  assign CAMLine_m_24_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_24_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_25_clock = clock;
  assign CAMLine_m_25_reset = reset;
  assign CAMLine_m_25_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_25_io_wi = io_waddr[25]; // @[cam.scala 144:31]
  assign CAMLine_m_25_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_25_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_26_clock = clock;
  assign CAMLine_m_26_reset = reset;
  assign CAMLine_m_26_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_26_io_wi = io_waddr[26]; // @[cam.scala 144:31]
  assign CAMLine_m_26_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_26_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_27_clock = clock;
  assign CAMLine_m_27_reset = reset;
  assign CAMLine_m_27_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_27_io_wi = io_waddr[27]; // @[cam.scala 144:31]
  assign CAMLine_m_27_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_27_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_28_clock = clock;
  assign CAMLine_m_28_reset = reset;
  assign CAMLine_m_28_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_28_io_wi = io_waddr[28]; // @[cam.scala 144:31]
  assign CAMLine_m_28_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_28_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_29_clock = clock;
  assign CAMLine_m_29_reset = reset;
  assign CAMLine_m_29_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_29_io_wi = io_waddr[29]; // @[cam.scala 144:31]
  assign CAMLine_m_29_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_29_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_30_clock = clock;
  assign CAMLine_m_30_reset = reset;
  assign CAMLine_m_30_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_30_io_wi = io_waddr[30]; // @[cam.scala 144:31]
  assign CAMLine_m_30_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_30_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_31_clock = clock;
  assign CAMLine_m_31_reset = reset;
  assign CAMLine_m_31_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_31_io_wi = io_waddr[31]; // @[cam.scala 144:31]
  assign CAMLine_m_31_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_31_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_32_clock = clock;
  assign CAMLine_m_32_reset = reset;
  assign CAMLine_m_32_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_32_io_wi = io_waddr[32]; // @[cam.scala 144:31]
  assign CAMLine_m_32_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_32_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_33_clock = clock;
  assign CAMLine_m_33_reset = reset;
  assign CAMLine_m_33_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_33_io_wi = io_waddr[33]; // @[cam.scala 144:31]
  assign CAMLine_m_33_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_33_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_34_clock = clock;
  assign CAMLine_m_34_reset = reset;
  assign CAMLine_m_34_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_34_io_wi = io_waddr[34]; // @[cam.scala 144:31]
  assign CAMLine_m_34_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_34_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_35_clock = clock;
  assign CAMLine_m_35_reset = reset;
  assign CAMLine_m_35_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_35_io_wi = io_waddr[35]; // @[cam.scala 144:31]
  assign CAMLine_m_35_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_35_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_36_clock = clock;
  assign CAMLine_m_36_reset = reset;
  assign CAMLine_m_36_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_36_io_wi = io_waddr[36]; // @[cam.scala 144:31]
  assign CAMLine_m_36_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_36_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_37_clock = clock;
  assign CAMLine_m_37_reset = reset;
  assign CAMLine_m_37_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_37_io_wi = io_waddr[37]; // @[cam.scala 144:31]
  assign CAMLine_m_37_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_37_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_38_clock = clock;
  assign CAMLine_m_38_reset = reset;
  assign CAMLine_m_38_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_38_io_wi = io_waddr[38]; // @[cam.scala 144:31]
  assign CAMLine_m_38_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_38_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_39_clock = clock;
  assign CAMLine_m_39_reset = reset;
  assign CAMLine_m_39_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_39_io_wi = io_waddr[39]; // @[cam.scala 144:31]
  assign CAMLine_m_39_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_39_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_40_clock = clock;
  assign CAMLine_m_40_reset = reset;
  assign CAMLine_m_40_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_40_io_wi = io_waddr[40]; // @[cam.scala 144:31]
  assign CAMLine_m_40_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_40_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_41_clock = clock;
  assign CAMLine_m_41_reset = reset;
  assign CAMLine_m_41_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_41_io_wi = io_waddr[41]; // @[cam.scala 144:31]
  assign CAMLine_m_41_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_41_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_42_clock = clock;
  assign CAMLine_m_42_reset = reset;
  assign CAMLine_m_42_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_42_io_wi = io_waddr[42]; // @[cam.scala 144:31]
  assign CAMLine_m_42_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_42_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_43_clock = clock;
  assign CAMLine_m_43_reset = reset;
  assign CAMLine_m_43_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_43_io_wi = io_waddr[43]; // @[cam.scala 144:31]
  assign CAMLine_m_43_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_43_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_44_clock = clock;
  assign CAMLine_m_44_reset = reset;
  assign CAMLine_m_44_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_44_io_wi = io_waddr[44]; // @[cam.scala 144:31]
  assign CAMLine_m_44_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_44_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_45_clock = clock;
  assign CAMLine_m_45_reset = reset;
  assign CAMLine_m_45_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_45_io_wi = io_waddr[45]; // @[cam.scala 144:31]
  assign CAMLine_m_45_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_45_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_46_clock = clock;
  assign CAMLine_m_46_reset = reset;
  assign CAMLine_m_46_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_46_io_wi = io_waddr[46]; // @[cam.scala 144:31]
  assign CAMLine_m_46_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_46_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_47_clock = clock;
  assign CAMLine_m_47_reset = reset;
  assign CAMLine_m_47_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_47_io_wi = io_waddr[47]; // @[cam.scala 144:31]
  assign CAMLine_m_47_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_47_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_48_clock = clock;
  assign CAMLine_m_48_reset = reset;
  assign CAMLine_m_48_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_48_io_wi = io_waddr[48]; // @[cam.scala 144:31]
  assign CAMLine_m_48_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_48_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_49_clock = clock;
  assign CAMLine_m_49_reset = reset;
  assign CAMLine_m_49_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_49_io_wi = io_waddr[49]; // @[cam.scala 144:31]
  assign CAMLine_m_49_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_49_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_50_clock = clock;
  assign CAMLine_m_50_reset = reset;
  assign CAMLine_m_50_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_50_io_wi = io_waddr[50]; // @[cam.scala 144:31]
  assign CAMLine_m_50_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_50_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_51_clock = clock;
  assign CAMLine_m_51_reset = reset;
  assign CAMLine_m_51_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_51_io_wi = io_waddr[51]; // @[cam.scala 144:31]
  assign CAMLine_m_51_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_51_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_52_clock = clock;
  assign CAMLine_m_52_reset = reset;
  assign CAMLine_m_52_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_52_io_wi = io_waddr[52]; // @[cam.scala 144:31]
  assign CAMLine_m_52_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_52_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_53_clock = clock;
  assign CAMLine_m_53_reset = reset;
  assign CAMLine_m_53_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_53_io_wi = io_waddr[53]; // @[cam.scala 144:31]
  assign CAMLine_m_53_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_53_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_54_clock = clock;
  assign CAMLine_m_54_reset = reset;
  assign CAMLine_m_54_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_54_io_wi = io_waddr[54]; // @[cam.scala 144:31]
  assign CAMLine_m_54_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_54_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_55_clock = clock;
  assign CAMLine_m_55_reset = reset;
  assign CAMLine_m_55_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_55_io_wi = io_waddr[55]; // @[cam.scala 144:31]
  assign CAMLine_m_55_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_55_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_56_clock = clock;
  assign CAMLine_m_56_reset = reset;
  assign CAMLine_m_56_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_56_io_wi = io_waddr[56]; // @[cam.scala 144:31]
  assign CAMLine_m_56_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_56_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_57_clock = clock;
  assign CAMLine_m_57_reset = reset;
  assign CAMLine_m_57_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_57_io_wi = io_waddr[57]; // @[cam.scala 144:31]
  assign CAMLine_m_57_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_57_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_58_clock = clock;
  assign CAMLine_m_58_reset = reset;
  assign CAMLine_m_58_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_58_io_wi = io_waddr[58]; // @[cam.scala 144:31]
  assign CAMLine_m_58_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_58_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_59_clock = clock;
  assign CAMLine_m_59_reset = reset;
  assign CAMLine_m_59_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_59_io_wi = io_waddr[59]; // @[cam.scala 144:31]
  assign CAMLine_m_59_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_59_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_60_clock = clock;
  assign CAMLine_m_60_reset = reset;
  assign CAMLine_m_60_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_60_io_wi = io_waddr[60]; // @[cam.scala 144:31]
  assign CAMLine_m_60_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_60_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_61_clock = clock;
  assign CAMLine_m_61_reset = reset;
  assign CAMLine_m_61_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_61_io_wi = io_waddr[61]; // @[cam.scala 144:31]
  assign CAMLine_m_61_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_61_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_62_clock = clock;
  assign CAMLine_m_62_reset = reset;
  assign CAMLine_m_62_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_62_io_wi = io_waddr[62]; // @[cam.scala 144:31]
  assign CAMLine_m_62_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_62_io_din = io_din; // @[cam.scala 146:21]
  assign CAMLine_m_63_clock = clock;
  assign CAMLine_m_63_reset = reset;
  assign CAMLine_m_63_io_we = io_we; // @[cam.scala 143:20]
  assign CAMLine_m_63_io_wi = io_waddr[63]; // @[cam.scala 144:31]
  assign CAMLine_m_63_io_key = io_key; // @[cam.scala 145:21]
  assign CAMLine_m_63_io_din = io_din; // @[cam.scala 146:21]
endmodule
