module RISCVCPUv2(
  input         clock,
  input         reset,
  input         io_rvfi_rst,
  input  [31:0] io_rvfi_insn_in_0,
  input  [31:0] io_rvfi_insn_in_1,
  input  [31:0] io_rvfi_insn_in_2,
  input  [31:0] io_rvfi_insn_in_3,
  input  [31:0] io_rvfi_insn_in_4,
  input  [31:0] io_rvfi_insn_in_5,
  input  [31:0] io_rvfi_insn_in_6,
  input  [31:0] io_rvfi_insn_in_7,
  input  [63:0] io_rvfi_reg_data_in_0,
  input  [63:0] io_rvfi_reg_data_in_1,
  input  [63:0] io_rvfi_reg_data_in_2,
  input  [63:0] io_rvfi_reg_data_in_3,
  input  [63:0] io_rvfi_reg_data_in_4,
  input  [63:0] io_rvfi_reg_data_in_5,
  input  [63:0] io_rvfi_reg_data_in_6,
  input  [63:0] io_rvfi_reg_data_in_7,
  input  [63:0] io_rvfi_reg_data_in_8,
  input  [63:0] io_rvfi_reg_data_in_9,
  input  [63:0] io_rvfi_reg_data_in_10,
  input  [63:0] io_rvfi_reg_data_in_11,
  input  [63:0] io_rvfi_reg_data_in_12,
  input  [63:0] io_rvfi_reg_data_in_13,
  input  [63:0] io_rvfi_reg_data_in_14,
  input  [63:0] io_rvfi_reg_data_in_15,
  input  [63:0] io_rvfi_reg_data_in_16,
  input  [63:0] io_rvfi_reg_data_in_17,
  input  [63:0] io_rvfi_reg_data_in_18,
  input  [63:0] io_rvfi_reg_data_in_19,
  input  [63:0] io_rvfi_reg_data_in_20,
  input  [63:0] io_rvfi_reg_data_in_21,
  input  [63:0] io_rvfi_reg_data_in_22,
  input  [63:0] io_rvfi_reg_data_in_23,
  input  [63:0] io_rvfi_reg_data_in_24,
  input  [63:0] io_rvfi_reg_data_in_25,
  input  [63:0] io_rvfi_reg_data_in_26,
  input  [63:0] io_rvfi_reg_data_in_27,
  input  [63:0] io_rvfi_reg_data_in_28,
  input  [63:0] io_rvfi_reg_data_in_29,
  input  [63:0] io_rvfi_reg_data_in_30,
  input  [63:0] io_rvfi_reg_data_in_31,
  input  [31:0] io_rvfi_mem_data_in_0,
  input  [31:0] io_rvfi_mem_data_in_1,
  input  [31:0] io_rvfi_mem_data_in_2,
  input  [31:0] io_rvfi_mem_data_in_3,
  input  [31:0] io_rvfi_mem_data_in_4,
  input  [31:0] io_rvfi_mem_data_in_5,
  input  [31:0] io_rvfi_mem_data_in_6,
  input  [31:0] io_rvfi_mem_data_in_7,
  input  [31:0] io_rvfi_mem_data_in_8,
  input  [31:0] io_rvfi_mem_data_in_9,
  input  [31:0] io_rvfi_mem_data_in_10,
  input  [31:0] io_rvfi_mem_data_in_11,
  input  [31:0] io_rvfi_mem_data_in_12,
  input  [31:0] io_rvfi_mem_data_in_13,
  input  [31:0] io_rvfi_mem_data_in_14,
  input  [31:0] io_rvfi_mem_data_in_15,
  input  [31:0] io_rvfi_mem_data_in_16,
  input  [31:0] io_rvfi_mem_data_in_17,
  input  [31:0] io_rvfi_mem_data_in_18,
  input  [31:0] io_rvfi_mem_data_in_19,
  input  [31:0] io_rvfi_mem_data_in_20,
  input  [31:0] io_rvfi_mem_data_in_21,
  input  [31:0] io_rvfi_mem_data_in_22,
  input  [31:0] io_rvfi_mem_data_in_23,
  input  [31:0] io_rvfi_mem_data_in_24,
  input  [31:0] io_rvfi_mem_data_in_25,
  input  [31:0] io_rvfi_mem_data_in_26,
  input  [31:0] io_rvfi_mem_data_in_27,
  input  [31:0] io_rvfi_mem_data_in_28,
  input  [31:0] io_rvfi_mem_data_in_29,
  input  [31:0] io_rvfi_mem_data_in_30,
  input  [31:0] io_rvfi_mem_data_in_31,
  input  [31:0] io_rvfi_mem_data_in_32,
  input  [31:0] io_rvfi_mem_data_in_33,
  input  [31:0] io_rvfi_mem_data_in_34,
  input  [31:0] io_rvfi_mem_data_in_35,
  input  [31:0] io_rvfi_mem_data_in_36,
  input  [31:0] io_rvfi_mem_data_in_37,
  input  [31:0] io_rvfi_mem_data_in_38,
  input  [31:0] io_rvfi_mem_data_in_39,
  input  [31:0] io_rvfi_mem_data_in_40,
  input  [31:0] io_rvfi_mem_data_in_41,
  input  [31:0] io_rvfi_mem_data_in_42,
  input  [31:0] io_rvfi_mem_data_in_43,
  input  [31:0] io_rvfi_mem_data_in_44,
  input  [31:0] io_rvfi_mem_data_in_45,
  input  [31:0] io_rvfi_mem_data_in_46,
  input  [31:0] io_rvfi_mem_data_in_47,
  input  [31:0] io_rvfi_mem_data_in_48,
  input  [31:0] io_rvfi_mem_data_in_49,
  input  [31:0] io_rvfi_mem_data_in_50,
  input  [31:0] io_rvfi_mem_data_in_51,
  input  [31:0] io_rvfi_mem_data_in_52,
  input  [31:0] io_rvfi_mem_data_in_53,
  input  [31:0] io_rvfi_mem_data_in_54,
  input  [31:0] io_rvfi_mem_data_in_55,
  input  [31:0] io_rvfi_mem_data_in_56,
  input  [31:0] io_rvfi_mem_data_in_57,
  input  [31:0] io_rvfi_mem_data_in_58,
  input  [31:0] io_rvfi_mem_data_in_59,
  input  [31:0] io_rvfi_mem_data_in_60,
  input  [31:0] io_rvfi_mem_data_in_61,
  input  [31:0] io_rvfi_mem_data_in_62,
  input  [31:0] io_rvfi_mem_data_in_63,
  input  [31:0] io_rvfi_mem_data_in_64,
  input  [31:0] io_rvfi_mem_data_in_65,
  input  [31:0] io_rvfi_mem_data_in_66,
  input  [31:0] io_rvfi_mem_data_in_67,
  input  [31:0] io_rvfi_mem_data_in_68,
  input  [31:0] io_rvfi_mem_data_in_69,
  input  [31:0] io_rvfi_mem_data_in_70,
  input  [31:0] io_rvfi_mem_data_in_71,
  input  [31:0] io_rvfi_mem_data_in_72,
  input  [31:0] io_rvfi_mem_data_in_73,
  input  [31:0] io_rvfi_mem_data_in_74,
  input  [31:0] io_rvfi_mem_data_in_75,
  input  [31:0] io_rvfi_mem_data_in_76,
  input  [31:0] io_rvfi_mem_data_in_77,
  input  [31:0] io_rvfi_mem_data_in_78,
  input  [31:0] io_rvfi_mem_data_in_79,
  input  [31:0] io_rvfi_mem_data_in_80,
  input  [31:0] io_rvfi_mem_data_in_81,
  input  [31:0] io_rvfi_mem_data_in_82,
  input  [31:0] io_rvfi_mem_data_in_83,
  input  [31:0] io_rvfi_mem_data_in_84,
  input  [31:0] io_rvfi_mem_data_in_85,
  input  [31:0] io_rvfi_mem_data_in_86,
  input  [31:0] io_rvfi_mem_data_in_87,
  input  [31:0] io_rvfi_mem_data_in_88,
  input  [31:0] io_rvfi_mem_data_in_89,
  input  [31:0] io_rvfi_mem_data_in_90,
  input  [31:0] io_rvfi_mem_data_in_91,
  input  [31:0] io_rvfi_mem_data_in_92,
  input  [31:0] io_rvfi_mem_data_in_93,
  input  [31:0] io_rvfi_mem_data_in_94,
  input  [31:0] io_rvfi_mem_data_in_95,
  input  [31:0] io_rvfi_mem_data_in_96,
  input  [31:0] io_rvfi_mem_data_in_97,
  input  [31:0] io_rvfi_mem_data_in_98,
  input  [31:0] io_rvfi_mem_data_in_99,
  input  [31:0] io_rvfi_mem_data_in_100,
  input  [31:0] io_rvfi_mem_data_in_101,
  input  [31:0] io_rvfi_mem_data_in_102,
  input  [31:0] io_rvfi_mem_data_in_103,
  input  [31:0] io_rvfi_mem_data_in_104,
  input  [31:0] io_rvfi_mem_data_in_105,
  input  [31:0] io_rvfi_mem_data_in_106,
  input  [31:0] io_rvfi_mem_data_in_107,
  input  [31:0] io_rvfi_mem_data_in_108,
  input  [31:0] io_rvfi_mem_data_in_109,
  input  [31:0] io_rvfi_mem_data_in_110,
  input  [31:0] io_rvfi_mem_data_in_111,
  input  [31:0] io_rvfi_mem_data_in_112,
  input  [31:0] io_rvfi_mem_data_in_113,
  input  [31:0] io_rvfi_mem_data_in_114,
  input  [31:0] io_rvfi_mem_data_in_115,
  input  [31:0] io_rvfi_mem_data_in_116,
  input  [31:0] io_rvfi_mem_data_in_117,
  input  [31:0] io_rvfi_mem_data_in_118,
  input  [31:0] io_rvfi_mem_data_in_119,
  input  [31:0] io_rvfi_mem_data_in_120,
  input  [31:0] io_rvfi_mem_data_in_121,
  input  [31:0] io_rvfi_mem_data_in_122,
  input  [31:0] io_rvfi_mem_data_in_123,
  input  [31:0] io_rvfi_mem_data_in_124,
  input  [31:0] io_rvfi_mem_data_in_125,
  input  [31:0] io_rvfi_mem_data_in_126,
  input  [31:0] io_rvfi_mem_data_in_127,
  input  [31:0] io_rvfi_mem_data_in_128,
  input  [31:0] io_rvfi_mem_data_in_129,
  input  [31:0] io_rvfi_mem_data_in_130,
  input  [31:0] io_rvfi_mem_data_in_131,
  input  [31:0] io_rvfi_mem_data_in_132,
  input  [31:0] io_rvfi_mem_data_in_133,
  input  [31:0] io_rvfi_mem_data_in_134,
  input  [31:0] io_rvfi_mem_data_in_135,
  input  [31:0] io_rvfi_mem_data_in_136,
  input  [31:0] io_rvfi_mem_data_in_137,
  input  [31:0] io_rvfi_mem_data_in_138,
  input  [31:0] io_rvfi_mem_data_in_139,
  input  [31:0] io_rvfi_mem_data_in_140,
  input  [31:0] io_rvfi_mem_data_in_141,
  input  [31:0] io_rvfi_mem_data_in_142,
  input  [31:0] io_rvfi_mem_data_in_143,
  input  [31:0] io_rvfi_mem_data_in_144,
  input  [31:0] io_rvfi_mem_data_in_145,
  input  [31:0] io_rvfi_mem_data_in_146,
  input  [31:0] io_rvfi_mem_data_in_147,
  input  [31:0] io_rvfi_mem_data_in_148,
  input  [31:0] io_rvfi_mem_data_in_149,
  input  [31:0] io_rvfi_mem_data_in_150,
  input  [31:0] io_rvfi_mem_data_in_151,
  input  [31:0] io_rvfi_mem_data_in_152,
  input  [31:0] io_rvfi_mem_data_in_153,
  input  [31:0] io_rvfi_mem_data_in_154,
  input  [31:0] io_rvfi_mem_data_in_155,
  input  [31:0] io_rvfi_mem_data_in_156,
  input  [31:0] io_rvfi_mem_data_in_157,
  input  [31:0] io_rvfi_mem_data_in_158,
  input  [31:0] io_rvfi_mem_data_in_159,
  input  [31:0] io_rvfi_mem_data_in_160,
  input  [31:0] io_rvfi_mem_data_in_161,
  input  [31:0] io_rvfi_mem_data_in_162,
  input  [31:0] io_rvfi_mem_data_in_163,
  input  [31:0] io_rvfi_mem_data_in_164,
  input  [31:0] io_rvfi_mem_data_in_165,
  input  [31:0] io_rvfi_mem_data_in_166,
  input  [31:0] io_rvfi_mem_data_in_167,
  input  [31:0] io_rvfi_mem_data_in_168,
  input  [31:0] io_rvfi_mem_data_in_169,
  input  [31:0] io_rvfi_mem_data_in_170,
  input  [31:0] io_rvfi_mem_data_in_171,
  input  [31:0] io_rvfi_mem_data_in_172,
  input  [31:0] io_rvfi_mem_data_in_173,
  input  [31:0] io_rvfi_mem_data_in_174,
  input  [31:0] io_rvfi_mem_data_in_175,
  input  [31:0] io_rvfi_mem_data_in_176,
  input  [31:0] io_rvfi_mem_data_in_177,
  input  [31:0] io_rvfi_mem_data_in_178,
  input  [31:0] io_rvfi_mem_data_in_179,
  input  [31:0] io_rvfi_mem_data_in_180,
  input  [31:0] io_rvfi_mem_data_in_181,
  input  [31:0] io_rvfi_mem_data_in_182,
  input  [31:0] io_rvfi_mem_data_in_183,
  input  [31:0] io_rvfi_mem_data_in_184,
  input  [31:0] io_rvfi_mem_data_in_185,
  input  [31:0] io_rvfi_mem_data_in_186,
  input  [31:0] io_rvfi_mem_data_in_187,
  input  [31:0] io_rvfi_mem_data_in_188,
  input  [31:0] io_rvfi_mem_data_in_189,
  input  [31:0] io_rvfi_mem_data_in_190,
  input  [31:0] io_rvfi_mem_data_in_191,
  input  [31:0] io_rvfi_mem_data_in_192,
  input  [31:0] io_rvfi_mem_data_in_193,
  input  [31:0] io_rvfi_mem_data_in_194,
  input  [31:0] io_rvfi_mem_data_in_195,
  input  [31:0] io_rvfi_mem_data_in_196,
  input  [31:0] io_rvfi_mem_data_in_197,
  input  [31:0] io_rvfi_mem_data_in_198,
  input  [31:0] io_rvfi_mem_data_in_199,
  input  [31:0] io_rvfi_mem_data_in_200,
  input  [31:0] io_rvfi_mem_data_in_201,
  input  [31:0] io_rvfi_mem_data_in_202,
  input  [31:0] io_rvfi_mem_data_in_203,
  input  [31:0] io_rvfi_mem_data_in_204,
  input  [31:0] io_rvfi_mem_data_in_205,
  input  [31:0] io_rvfi_mem_data_in_206,
  input  [31:0] io_rvfi_mem_data_in_207,
  input  [31:0] io_rvfi_mem_data_in_208,
  input  [31:0] io_rvfi_mem_data_in_209,
  input  [31:0] io_rvfi_mem_data_in_210,
  input  [31:0] io_rvfi_mem_data_in_211,
  input  [31:0] io_rvfi_mem_data_in_212,
  input  [31:0] io_rvfi_mem_data_in_213,
  input  [31:0] io_rvfi_mem_data_in_214,
  input  [31:0] io_rvfi_mem_data_in_215,
  input  [31:0] io_rvfi_mem_data_in_216,
  input  [31:0] io_rvfi_mem_data_in_217,
  input  [31:0] io_rvfi_mem_data_in_218,
  input  [31:0] io_rvfi_mem_data_in_219,
  input  [31:0] io_rvfi_mem_data_in_220,
  input  [31:0] io_rvfi_mem_data_in_221,
  input  [31:0] io_rvfi_mem_data_in_222,
  input  [31:0] io_rvfi_mem_data_in_223,
  input  [31:0] io_rvfi_mem_data_in_224,
  input  [31:0] io_rvfi_mem_data_in_225,
  input  [31:0] io_rvfi_mem_data_in_226,
  input  [31:0] io_rvfi_mem_data_in_227,
  input  [31:0] io_rvfi_mem_data_in_228,
  input  [31:0] io_rvfi_mem_data_in_229,
  input  [31:0] io_rvfi_mem_data_in_230,
  input  [31:0] io_rvfi_mem_data_in_231,
  input  [31:0] io_rvfi_mem_data_in_232,
  input  [31:0] io_rvfi_mem_data_in_233,
  input  [31:0] io_rvfi_mem_data_in_234,
  input  [31:0] io_rvfi_mem_data_in_235,
  input  [31:0] io_rvfi_mem_data_in_236,
  input  [31:0] io_rvfi_mem_data_in_237,
  input  [31:0] io_rvfi_mem_data_in_238,
  input  [31:0] io_rvfi_mem_data_in_239,
  input  [31:0] io_rvfi_mem_data_in_240,
  input  [31:0] io_rvfi_mem_data_in_241,
  input  [31:0] io_rvfi_mem_data_in_242,
  input  [31:0] io_rvfi_mem_data_in_243,
  input  [31:0] io_rvfi_mem_data_in_244,
  input  [31:0] io_rvfi_mem_data_in_245,
  input  [31:0] io_rvfi_mem_data_in_246,
  input  [31:0] io_rvfi_mem_data_in_247,
  input  [31:0] io_rvfi_mem_data_in_248,
  input  [31:0] io_rvfi_mem_data_in_249,
  input  [31:0] io_rvfi_mem_data_in_250,
  input  [31:0] io_rvfi_mem_data_in_251,
  input  [31:0] io_rvfi_mem_data_in_252,
  input  [31:0] io_rvfi_mem_data_in_253,
  input  [31:0] io_rvfi_mem_data_in_254,
  input  [31:0] io_rvfi_mem_data_in_255,
  input  [31:0] io_rvfi_mem_data_in_256,
  input  [31:0] io_rvfi_mem_data_in_257,
  input  [31:0] io_rvfi_mem_data_in_258,
  input  [31:0] io_rvfi_mem_data_in_259,
  input  [31:0] io_rvfi_mem_data_in_260,
  input  [31:0] io_rvfi_mem_data_in_261,
  input  [31:0] io_rvfi_mem_data_in_262,
  input  [31:0] io_rvfi_mem_data_in_263,
  input  [31:0] io_rvfi_mem_data_in_264,
  input  [31:0] io_rvfi_mem_data_in_265,
  input  [31:0] io_rvfi_mem_data_in_266,
  input  [31:0] io_rvfi_mem_data_in_267,
  input  [31:0] io_rvfi_mem_data_in_268,
  input  [31:0] io_rvfi_mem_data_in_269,
  input  [31:0] io_rvfi_mem_data_in_270,
  input  [31:0] io_rvfi_mem_data_in_271,
  input  [31:0] io_rvfi_mem_data_in_272,
  input  [31:0] io_rvfi_mem_data_in_273,
  input  [31:0] io_rvfi_mem_data_in_274,
  input  [31:0] io_rvfi_mem_data_in_275,
  input  [31:0] io_rvfi_mem_data_in_276,
  input  [31:0] io_rvfi_mem_data_in_277,
  input  [31:0] io_rvfi_mem_data_in_278,
  input  [31:0] io_rvfi_mem_data_in_279,
  input  [31:0] io_rvfi_mem_data_in_280,
  input  [31:0] io_rvfi_mem_data_in_281,
  input  [31:0] io_rvfi_mem_data_in_282,
  input  [31:0] io_rvfi_mem_data_in_283,
  input  [31:0] io_rvfi_mem_data_in_284,
  input  [31:0] io_rvfi_mem_data_in_285,
  input  [31:0] io_rvfi_mem_data_in_286,
  input  [31:0] io_rvfi_mem_data_in_287,
  input  [31:0] io_rvfi_mem_data_in_288,
  input  [31:0] io_rvfi_mem_data_in_289,
  input  [31:0] io_rvfi_mem_data_in_290,
  input  [31:0] io_rvfi_mem_data_in_291,
  input  [31:0] io_rvfi_mem_data_in_292,
  input  [31:0] io_rvfi_mem_data_in_293,
  input  [31:0] io_rvfi_mem_data_in_294,
  input  [31:0] io_rvfi_mem_data_in_295,
  input  [31:0] io_rvfi_mem_data_in_296,
  input  [31:0] io_rvfi_mem_data_in_297,
  input  [31:0] io_rvfi_mem_data_in_298,
  input  [31:0] io_rvfi_mem_data_in_299,
  input  [31:0] io_rvfi_mem_data_in_300,
  input  [31:0] io_rvfi_mem_data_in_301,
  input  [31:0] io_rvfi_mem_data_in_302,
  input  [31:0] io_rvfi_mem_data_in_303,
  input  [31:0] io_rvfi_mem_data_in_304,
  input  [31:0] io_rvfi_mem_data_in_305,
  input  [31:0] io_rvfi_mem_data_in_306,
  input  [31:0] io_rvfi_mem_data_in_307,
  input  [31:0] io_rvfi_mem_data_in_308,
  input  [31:0] io_rvfi_mem_data_in_309,
  input  [31:0] io_rvfi_mem_data_in_310,
  input  [31:0] io_rvfi_mem_data_in_311,
  input  [31:0] io_rvfi_mem_data_in_312,
  input  [31:0] io_rvfi_mem_data_in_313,
  input  [31:0] io_rvfi_mem_data_in_314,
  input  [31:0] io_rvfi_mem_data_in_315,
  input  [31:0] io_rvfi_mem_data_in_316,
  input  [31:0] io_rvfi_mem_data_in_317,
  input  [31:0] io_rvfi_mem_data_in_318,
  input  [31:0] io_rvfi_mem_data_in_319,
  input  [31:0] io_rvfi_mem_data_in_320,
  input  [31:0] io_rvfi_mem_data_in_321,
  input  [31:0] io_rvfi_mem_data_in_322,
  input  [31:0] io_rvfi_mem_data_in_323,
  input  [31:0] io_rvfi_mem_data_in_324,
  input  [31:0] io_rvfi_mem_data_in_325,
  input  [31:0] io_rvfi_mem_data_in_326,
  input  [31:0] io_rvfi_mem_data_in_327,
  input  [31:0] io_rvfi_mem_data_in_328,
  input  [31:0] io_rvfi_mem_data_in_329,
  input  [31:0] io_rvfi_mem_data_in_330,
  input  [31:0] io_rvfi_mem_data_in_331,
  input  [31:0] io_rvfi_mem_data_in_332,
  input  [31:0] io_rvfi_mem_data_in_333,
  input  [31:0] io_rvfi_mem_data_in_334,
  input  [31:0] io_rvfi_mem_data_in_335,
  input  [31:0] io_rvfi_mem_data_in_336,
  input  [31:0] io_rvfi_mem_data_in_337,
  input  [31:0] io_rvfi_mem_data_in_338,
  input  [31:0] io_rvfi_mem_data_in_339,
  input  [31:0] io_rvfi_mem_data_in_340,
  input  [31:0] io_rvfi_mem_data_in_341,
  input  [31:0] io_rvfi_mem_data_in_342,
  input  [31:0] io_rvfi_mem_data_in_343,
  input  [31:0] io_rvfi_mem_data_in_344,
  input  [31:0] io_rvfi_mem_data_in_345,
  input  [31:0] io_rvfi_mem_data_in_346,
  input  [31:0] io_rvfi_mem_data_in_347,
  input  [31:0] io_rvfi_mem_data_in_348,
  input  [31:0] io_rvfi_mem_data_in_349,
  input  [31:0] io_rvfi_mem_data_in_350,
  input  [31:0] io_rvfi_mem_data_in_351,
  input  [31:0] io_rvfi_mem_data_in_352,
  input  [31:0] io_rvfi_mem_data_in_353,
  input  [31:0] io_rvfi_mem_data_in_354,
  input  [31:0] io_rvfi_mem_data_in_355,
  input  [31:0] io_rvfi_mem_data_in_356,
  input  [31:0] io_rvfi_mem_data_in_357,
  input  [31:0] io_rvfi_mem_data_in_358,
  input  [31:0] io_rvfi_mem_data_in_359,
  input  [31:0] io_rvfi_mem_data_in_360,
  input  [31:0] io_rvfi_mem_data_in_361,
  input  [31:0] io_rvfi_mem_data_in_362,
  input  [31:0] io_rvfi_mem_data_in_363,
  input  [31:0] io_rvfi_mem_data_in_364,
  input  [31:0] io_rvfi_mem_data_in_365,
  input  [31:0] io_rvfi_mem_data_in_366,
  input  [31:0] io_rvfi_mem_data_in_367,
  input  [31:0] io_rvfi_mem_data_in_368,
  input  [31:0] io_rvfi_mem_data_in_369,
  input  [31:0] io_rvfi_mem_data_in_370,
  input  [31:0] io_rvfi_mem_data_in_371,
  input  [31:0] io_rvfi_mem_data_in_372,
  input  [31:0] io_rvfi_mem_data_in_373,
  input  [31:0] io_rvfi_mem_data_in_374,
  input  [31:0] io_rvfi_mem_data_in_375,
  input  [31:0] io_rvfi_mem_data_in_376,
  input  [31:0] io_rvfi_mem_data_in_377,
  input  [31:0] io_rvfi_mem_data_in_378,
  input  [31:0] io_rvfi_mem_data_in_379,
  input  [31:0] io_rvfi_mem_data_in_380,
  input  [31:0] io_rvfi_mem_data_in_381,
  input  [31:0] io_rvfi_mem_data_in_382,
  input  [31:0] io_rvfi_mem_data_in_383,
  input  [31:0] io_rvfi_mem_data_in_384,
  input  [31:0] io_rvfi_mem_data_in_385,
  input  [31:0] io_rvfi_mem_data_in_386,
  input  [31:0] io_rvfi_mem_data_in_387,
  input  [31:0] io_rvfi_mem_data_in_388,
  input  [31:0] io_rvfi_mem_data_in_389,
  input  [31:0] io_rvfi_mem_data_in_390,
  input  [31:0] io_rvfi_mem_data_in_391,
  input  [31:0] io_rvfi_mem_data_in_392,
  input  [31:0] io_rvfi_mem_data_in_393,
  input  [31:0] io_rvfi_mem_data_in_394,
  input  [31:0] io_rvfi_mem_data_in_395,
  input  [31:0] io_rvfi_mem_data_in_396,
  input  [31:0] io_rvfi_mem_data_in_397,
  input  [31:0] io_rvfi_mem_data_in_398,
  input  [31:0] io_rvfi_mem_data_in_399,
  input  [31:0] io_rvfi_mem_data_in_400,
  input  [31:0] io_rvfi_mem_data_in_401,
  input  [31:0] io_rvfi_mem_data_in_402,
  input  [31:0] io_rvfi_mem_data_in_403,
  input  [31:0] io_rvfi_mem_data_in_404,
  input  [31:0] io_rvfi_mem_data_in_405,
  input  [31:0] io_rvfi_mem_data_in_406,
  input  [31:0] io_rvfi_mem_data_in_407,
  input  [31:0] io_rvfi_mem_data_in_408,
  input  [31:0] io_rvfi_mem_data_in_409,
  input  [31:0] io_rvfi_mem_data_in_410,
  input  [31:0] io_rvfi_mem_data_in_411,
  input  [31:0] io_rvfi_mem_data_in_412,
  input  [31:0] io_rvfi_mem_data_in_413,
  input  [31:0] io_rvfi_mem_data_in_414,
  input  [31:0] io_rvfi_mem_data_in_415,
  input  [31:0] io_rvfi_mem_data_in_416,
  input  [31:0] io_rvfi_mem_data_in_417,
  input  [31:0] io_rvfi_mem_data_in_418,
  input  [31:0] io_rvfi_mem_data_in_419,
  input  [31:0] io_rvfi_mem_data_in_420,
  input  [31:0] io_rvfi_mem_data_in_421,
  input  [31:0] io_rvfi_mem_data_in_422,
  input  [31:0] io_rvfi_mem_data_in_423,
  input  [31:0] io_rvfi_mem_data_in_424,
  input  [31:0] io_rvfi_mem_data_in_425,
  input  [31:0] io_rvfi_mem_data_in_426,
  input  [31:0] io_rvfi_mem_data_in_427,
  input  [31:0] io_rvfi_mem_data_in_428,
  input  [31:0] io_rvfi_mem_data_in_429,
  input  [31:0] io_rvfi_mem_data_in_430,
  input  [31:0] io_rvfi_mem_data_in_431,
  input  [31:0] io_rvfi_mem_data_in_432,
  input  [31:0] io_rvfi_mem_data_in_433,
  input  [31:0] io_rvfi_mem_data_in_434,
  input  [31:0] io_rvfi_mem_data_in_435,
  input  [31:0] io_rvfi_mem_data_in_436,
  input  [31:0] io_rvfi_mem_data_in_437,
  input  [31:0] io_rvfi_mem_data_in_438,
  input  [31:0] io_rvfi_mem_data_in_439,
  input  [31:0] io_rvfi_mem_data_in_440,
  input  [31:0] io_rvfi_mem_data_in_441,
  input  [31:0] io_rvfi_mem_data_in_442,
  input  [31:0] io_rvfi_mem_data_in_443,
  input  [31:0] io_rvfi_mem_data_in_444,
  input  [31:0] io_rvfi_mem_data_in_445,
  input  [31:0] io_rvfi_mem_data_in_446,
  input  [31:0] io_rvfi_mem_data_in_447,
  input  [31:0] io_rvfi_mem_data_in_448,
  input  [31:0] io_rvfi_mem_data_in_449,
  input  [31:0] io_rvfi_mem_data_in_450,
  input  [31:0] io_rvfi_mem_data_in_451,
  input  [31:0] io_rvfi_mem_data_in_452,
  input  [31:0] io_rvfi_mem_data_in_453,
  input  [31:0] io_rvfi_mem_data_in_454,
  input  [31:0] io_rvfi_mem_data_in_455,
  input  [31:0] io_rvfi_mem_data_in_456,
  input  [31:0] io_rvfi_mem_data_in_457,
  input  [31:0] io_rvfi_mem_data_in_458,
  input  [31:0] io_rvfi_mem_data_in_459,
  input  [31:0] io_rvfi_mem_data_in_460,
  input  [31:0] io_rvfi_mem_data_in_461,
  input  [31:0] io_rvfi_mem_data_in_462,
  input  [31:0] io_rvfi_mem_data_in_463,
  input  [31:0] io_rvfi_mem_data_in_464,
  input  [31:0] io_rvfi_mem_data_in_465,
  input  [31:0] io_rvfi_mem_data_in_466,
  input  [31:0] io_rvfi_mem_data_in_467,
  input  [31:0] io_rvfi_mem_data_in_468,
  input  [31:0] io_rvfi_mem_data_in_469,
  input  [31:0] io_rvfi_mem_data_in_470,
  input  [31:0] io_rvfi_mem_data_in_471,
  input  [31:0] io_rvfi_mem_data_in_472,
  input  [31:0] io_rvfi_mem_data_in_473,
  input  [31:0] io_rvfi_mem_data_in_474,
  input  [31:0] io_rvfi_mem_data_in_475,
  input  [31:0] io_rvfi_mem_data_in_476,
  input  [31:0] io_rvfi_mem_data_in_477,
  input  [31:0] io_rvfi_mem_data_in_478,
  input  [31:0] io_rvfi_mem_data_in_479,
  input  [31:0] io_rvfi_mem_data_in_480,
  input  [31:0] io_rvfi_mem_data_in_481,
  input  [31:0] io_rvfi_mem_data_in_482,
  input  [31:0] io_rvfi_mem_data_in_483,
  input  [31:0] io_rvfi_mem_data_in_484,
  input  [31:0] io_rvfi_mem_data_in_485,
  input  [31:0] io_rvfi_mem_data_in_486,
  input  [31:0] io_rvfi_mem_data_in_487,
  input  [31:0] io_rvfi_mem_data_in_488,
  input  [31:0] io_rvfi_mem_data_in_489,
  input  [31:0] io_rvfi_mem_data_in_490,
  input  [31:0] io_rvfi_mem_data_in_491,
  input  [31:0] io_rvfi_mem_data_in_492,
  input  [31:0] io_rvfi_mem_data_in_493,
  input  [31:0] io_rvfi_mem_data_in_494,
  input  [31:0] io_rvfi_mem_data_in_495,
  input  [31:0] io_rvfi_mem_data_in_496,
  input  [31:0] io_rvfi_mem_data_in_497,
  input  [31:0] io_rvfi_mem_data_in_498,
  input  [31:0] io_rvfi_mem_data_in_499,
  input  [31:0] io_rvfi_mem_data_in_500,
  input  [31:0] io_rvfi_mem_data_in_501,
  input  [31:0] io_rvfi_mem_data_in_502,
  input  [31:0] io_rvfi_mem_data_in_503,
  input  [31:0] io_rvfi_mem_data_in_504,
  input  [31:0] io_rvfi_mem_data_in_505,
  input  [31:0] io_rvfi_mem_data_in_506,
  input  [31:0] io_rvfi_mem_data_in_507,
  input  [31:0] io_rvfi_mem_data_in_508,
  input  [31:0] io_rvfi_mem_data_in_509,
  input  [31:0] io_rvfi_mem_data_in_510,
  input  [31:0] io_rvfi_mem_data_in_511,
  input  [31:0] io_rvfi_mem_data_in_512,
  input  [31:0] io_rvfi_mem_data_in_513,
  input  [31:0] io_rvfi_mem_data_in_514,
  input  [31:0] io_rvfi_mem_data_in_515,
  input  [31:0] io_rvfi_mem_data_in_516,
  input  [31:0] io_rvfi_mem_data_in_517,
  input  [31:0] io_rvfi_mem_data_in_518,
  input  [31:0] io_rvfi_mem_data_in_519,
  input  [31:0] io_rvfi_mem_data_in_520,
  input  [31:0] io_rvfi_mem_data_in_521,
  input  [31:0] io_rvfi_mem_data_in_522,
  input  [31:0] io_rvfi_mem_data_in_523,
  input  [31:0] io_rvfi_mem_data_in_524,
  input  [31:0] io_rvfi_mem_data_in_525,
  input  [31:0] io_rvfi_mem_data_in_526,
  input  [31:0] io_rvfi_mem_data_in_527,
  input  [31:0] io_rvfi_mem_data_in_528,
  input  [31:0] io_rvfi_mem_data_in_529,
  input  [31:0] io_rvfi_mem_data_in_530,
  input  [31:0] io_rvfi_mem_data_in_531,
  input  [31:0] io_rvfi_mem_data_in_532,
  input  [31:0] io_rvfi_mem_data_in_533,
  input  [31:0] io_rvfi_mem_data_in_534,
  input  [31:0] io_rvfi_mem_data_in_535,
  input  [31:0] io_rvfi_mem_data_in_536,
  input  [31:0] io_rvfi_mem_data_in_537,
  input  [31:0] io_rvfi_mem_data_in_538,
  input  [31:0] io_rvfi_mem_data_in_539,
  input  [31:0] io_rvfi_mem_data_in_540,
  input  [31:0] io_rvfi_mem_data_in_541,
  input  [31:0] io_rvfi_mem_data_in_542,
  input  [31:0] io_rvfi_mem_data_in_543,
  input  [31:0] io_rvfi_mem_data_in_544,
  input  [31:0] io_rvfi_mem_data_in_545,
  input  [31:0] io_rvfi_mem_data_in_546,
  input  [31:0] io_rvfi_mem_data_in_547,
  input  [31:0] io_rvfi_mem_data_in_548,
  input  [31:0] io_rvfi_mem_data_in_549,
  input  [31:0] io_rvfi_mem_data_in_550,
  input  [31:0] io_rvfi_mem_data_in_551,
  input  [31:0] io_rvfi_mem_data_in_552,
  input  [31:0] io_rvfi_mem_data_in_553,
  input  [31:0] io_rvfi_mem_data_in_554,
  input  [31:0] io_rvfi_mem_data_in_555,
  input  [31:0] io_rvfi_mem_data_in_556,
  input  [31:0] io_rvfi_mem_data_in_557,
  input  [31:0] io_rvfi_mem_data_in_558,
  input  [31:0] io_rvfi_mem_data_in_559,
  input  [31:0] io_rvfi_mem_data_in_560,
  input  [31:0] io_rvfi_mem_data_in_561,
  input  [31:0] io_rvfi_mem_data_in_562,
  input  [31:0] io_rvfi_mem_data_in_563,
  input  [31:0] io_rvfi_mem_data_in_564,
  input  [31:0] io_rvfi_mem_data_in_565,
  input  [31:0] io_rvfi_mem_data_in_566,
  input  [31:0] io_rvfi_mem_data_in_567,
  input  [31:0] io_rvfi_mem_data_in_568,
  input  [31:0] io_rvfi_mem_data_in_569,
  input  [31:0] io_rvfi_mem_data_in_570,
  input  [31:0] io_rvfi_mem_data_in_571,
  input  [31:0] io_rvfi_mem_data_in_572,
  input  [31:0] io_rvfi_mem_data_in_573,
  input  [31:0] io_rvfi_mem_data_in_574,
  input  [31:0] io_rvfi_mem_data_in_575,
  input  [31:0] io_rvfi_mem_data_in_576,
  input  [31:0] io_rvfi_mem_data_in_577,
  input  [31:0] io_rvfi_mem_data_in_578,
  input  [31:0] io_rvfi_mem_data_in_579,
  input  [31:0] io_rvfi_mem_data_in_580,
  input  [31:0] io_rvfi_mem_data_in_581,
  input  [31:0] io_rvfi_mem_data_in_582,
  input  [31:0] io_rvfi_mem_data_in_583,
  input  [31:0] io_rvfi_mem_data_in_584,
  input  [31:0] io_rvfi_mem_data_in_585,
  input  [31:0] io_rvfi_mem_data_in_586,
  input  [31:0] io_rvfi_mem_data_in_587,
  input  [31:0] io_rvfi_mem_data_in_588,
  input  [31:0] io_rvfi_mem_data_in_589,
  input  [31:0] io_rvfi_mem_data_in_590,
  input  [31:0] io_rvfi_mem_data_in_591,
  input  [31:0] io_rvfi_mem_data_in_592,
  input  [31:0] io_rvfi_mem_data_in_593,
  input  [31:0] io_rvfi_mem_data_in_594,
  input  [31:0] io_rvfi_mem_data_in_595,
  input  [31:0] io_rvfi_mem_data_in_596,
  input  [31:0] io_rvfi_mem_data_in_597,
  input  [31:0] io_rvfi_mem_data_in_598,
  input  [31:0] io_rvfi_mem_data_in_599,
  input  [31:0] io_rvfi_mem_data_in_600,
  input  [31:0] io_rvfi_mem_data_in_601,
  input  [31:0] io_rvfi_mem_data_in_602,
  input  [31:0] io_rvfi_mem_data_in_603,
  input  [31:0] io_rvfi_mem_data_in_604,
  input  [31:0] io_rvfi_mem_data_in_605,
  input  [31:0] io_rvfi_mem_data_in_606,
  input  [31:0] io_rvfi_mem_data_in_607,
  input  [31:0] io_rvfi_mem_data_in_608,
  input  [31:0] io_rvfi_mem_data_in_609,
  input  [31:0] io_rvfi_mem_data_in_610,
  input  [31:0] io_rvfi_mem_data_in_611,
  input  [31:0] io_rvfi_mem_data_in_612,
  input  [31:0] io_rvfi_mem_data_in_613,
  input  [31:0] io_rvfi_mem_data_in_614,
  input  [31:0] io_rvfi_mem_data_in_615,
  input  [31:0] io_rvfi_mem_data_in_616,
  input  [31:0] io_rvfi_mem_data_in_617,
  input  [31:0] io_rvfi_mem_data_in_618,
  input  [31:0] io_rvfi_mem_data_in_619,
  input  [31:0] io_rvfi_mem_data_in_620,
  input  [31:0] io_rvfi_mem_data_in_621,
  input  [31:0] io_rvfi_mem_data_in_622,
  input  [31:0] io_rvfi_mem_data_in_623,
  input  [31:0] io_rvfi_mem_data_in_624,
  input  [31:0] io_rvfi_mem_data_in_625,
  input  [31:0] io_rvfi_mem_data_in_626,
  input  [31:0] io_rvfi_mem_data_in_627,
  input  [31:0] io_rvfi_mem_data_in_628,
  input  [31:0] io_rvfi_mem_data_in_629,
  input  [31:0] io_rvfi_mem_data_in_630,
  input  [31:0] io_rvfi_mem_data_in_631,
  input  [31:0] io_rvfi_mem_data_in_632,
  input  [31:0] io_rvfi_mem_data_in_633,
  input  [31:0] io_rvfi_mem_data_in_634,
  input  [31:0] io_rvfi_mem_data_in_635,
  input  [31:0] io_rvfi_mem_data_in_636,
  input  [31:0] io_rvfi_mem_data_in_637,
  input  [31:0] io_rvfi_mem_data_in_638,
  input  [31:0] io_rvfi_mem_data_in_639,
  input  [31:0] io_rvfi_mem_data_in_640,
  input  [31:0] io_rvfi_mem_data_in_641,
  input  [31:0] io_rvfi_mem_data_in_642,
  input  [31:0] io_rvfi_mem_data_in_643,
  input  [31:0] io_rvfi_mem_data_in_644,
  input  [31:0] io_rvfi_mem_data_in_645,
  input  [31:0] io_rvfi_mem_data_in_646,
  input  [31:0] io_rvfi_mem_data_in_647,
  input  [31:0] io_rvfi_mem_data_in_648,
  input  [31:0] io_rvfi_mem_data_in_649,
  input  [31:0] io_rvfi_mem_data_in_650,
  input  [31:0] io_rvfi_mem_data_in_651,
  input  [31:0] io_rvfi_mem_data_in_652,
  input  [31:0] io_rvfi_mem_data_in_653,
  input  [31:0] io_rvfi_mem_data_in_654,
  input  [31:0] io_rvfi_mem_data_in_655,
  input  [31:0] io_rvfi_mem_data_in_656,
  input  [31:0] io_rvfi_mem_data_in_657,
  input  [31:0] io_rvfi_mem_data_in_658,
  input  [31:0] io_rvfi_mem_data_in_659,
  input  [31:0] io_rvfi_mem_data_in_660,
  input  [31:0] io_rvfi_mem_data_in_661,
  input  [31:0] io_rvfi_mem_data_in_662,
  input  [31:0] io_rvfi_mem_data_in_663,
  input  [31:0] io_rvfi_mem_data_in_664,
  input  [31:0] io_rvfi_mem_data_in_665,
  input  [31:0] io_rvfi_mem_data_in_666,
  input  [31:0] io_rvfi_mem_data_in_667,
  input  [31:0] io_rvfi_mem_data_in_668,
  input  [31:0] io_rvfi_mem_data_in_669,
  input  [31:0] io_rvfi_mem_data_in_670,
  input  [31:0] io_rvfi_mem_data_in_671,
  input  [31:0] io_rvfi_mem_data_in_672,
  input  [31:0] io_rvfi_mem_data_in_673,
  input  [31:0] io_rvfi_mem_data_in_674,
  input  [31:0] io_rvfi_mem_data_in_675,
  input  [31:0] io_rvfi_mem_data_in_676,
  input  [31:0] io_rvfi_mem_data_in_677,
  input  [31:0] io_rvfi_mem_data_in_678,
  input  [31:0] io_rvfi_mem_data_in_679,
  input  [31:0] io_rvfi_mem_data_in_680,
  input  [31:0] io_rvfi_mem_data_in_681,
  input  [31:0] io_rvfi_mem_data_in_682,
  input  [31:0] io_rvfi_mem_data_in_683,
  input  [31:0] io_rvfi_mem_data_in_684,
  input  [31:0] io_rvfi_mem_data_in_685,
  input  [31:0] io_rvfi_mem_data_in_686,
  input  [31:0] io_rvfi_mem_data_in_687,
  input  [31:0] io_rvfi_mem_data_in_688,
  input  [31:0] io_rvfi_mem_data_in_689,
  input  [31:0] io_rvfi_mem_data_in_690,
  input  [31:0] io_rvfi_mem_data_in_691,
  input  [31:0] io_rvfi_mem_data_in_692,
  input  [31:0] io_rvfi_mem_data_in_693,
  input  [31:0] io_rvfi_mem_data_in_694,
  input  [31:0] io_rvfi_mem_data_in_695,
  input  [31:0] io_rvfi_mem_data_in_696,
  input  [31:0] io_rvfi_mem_data_in_697,
  input  [31:0] io_rvfi_mem_data_in_698,
  input  [31:0] io_rvfi_mem_data_in_699,
  input  [31:0] io_rvfi_mem_data_in_700,
  input  [31:0] io_rvfi_mem_data_in_701,
  input  [31:0] io_rvfi_mem_data_in_702,
  input  [31:0] io_rvfi_mem_data_in_703,
  input  [31:0] io_rvfi_mem_data_in_704,
  input  [31:0] io_rvfi_mem_data_in_705,
  input  [31:0] io_rvfi_mem_data_in_706,
  input  [31:0] io_rvfi_mem_data_in_707,
  input  [31:0] io_rvfi_mem_data_in_708,
  input  [31:0] io_rvfi_mem_data_in_709,
  input  [31:0] io_rvfi_mem_data_in_710,
  input  [31:0] io_rvfi_mem_data_in_711,
  input  [31:0] io_rvfi_mem_data_in_712,
  input  [31:0] io_rvfi_mem_data_in_713,
  input  [31:0] io_rvfi_mem_data_in_714,
  input  [31:0] io_rvfi_mem_data_in_715,
  input  [31:0] io_rvfi_mem_data_in_716,
  input  [31:0] io_rvfi_mem_data_in_717,
  input  [31:0] io_rvfi_mem_data_in_718,
  input  [31:0] io_rvfi_mem_data_in_719,
  input  [31:0] io_rvfi_mem_data_in_720,
  input  [31:0] io_rvfi_mem_data_in_721,
  input  [31:0] io_rvfi_mem_data_in_722,
  input  [31:0] io_rvfi_mem_data_in_723,
  input  [31:0] io_rvfi_mem_data_in_724,
  input  [31:0] io_rvfi_mem_data_in_725,
  input  [31:0] io_rvfi_mem_data_in_726,
  input  [31:0] io_rvfi_mem_data_in_727,
  input  [31:0] io_rvfi_mem_data_in_728,
  input  [31:0] io_rvfi_mem_data_in_729,
  input  [31:0] io_rvfi_mem_data_in_730,
  input  [31:0] io_rvfi_mem_data_in_731,
  input  [31:0] io_rvfi_mem_data_in_732,
  input  [31:0] io_rvfi_mem_data_in_733,
  input  [31:0] io_rvfi_mem_data_in_734,
  input  [31:0] io_rvfi_mem_data_in_735,
  input  [31:0] io_rvfi_mem_data_in_736,
  input  [31:0] io_rvfi_mem_data_in_737,
  input  [31:0] io_rvfi_mem_data_in_738,
  input  [31:0] io_rvfi_mem_data_in_739,
  input  [31:0] io_rvfi_mem_data_in_740,
  input  [31:0] io_rvfi_mem_data_in_741,
  input  [31:0] io_rvfi_mem_data_in_742,
  input  [31:0] io_rvfi_mem_data_in_743,
  input  [31:0] io_rvfi_mem_data_in_744,
  input  [31:0] io_rvfi_mem_data_in_745,
  input  [31:0] io_rvfi_mem_data_in_746,
  input  [31:0] io_rvfi_mem_data_in_747,
  input  [31:0] io_rvfi_mem_data_in_748,
  input  [31:0] io_rvfi_mem_data_in_749,
  input  [31:0] io_rvfi_mem_data_in_750,
  input  [31:0] io_rvfi_mem_data_in_751,
  input  [31:0] io_rvfi_mem_data_in_752,
  input  [31:0] io_rvfi_mem_data_in_753,
  input  [31:0] io_rvfi_mem_data_in_754,
  input  [31:0] io_rvfi_mem_data_in_755,
  input  [31:0] io_rvfi_mem_data_in_756,
  input  [31:0] io_rvfi_mem_data_in_757,
  input  [31:0] io_rvfi_mem_data_in_758,
  input  [31:0] io_rvfi_mem_data_in_759,
  input  [31:0] io_rvfi_mem_data_in_760,
  input  [31:0] io_rvfi_mem_data_in_761,
  input  [31:0] io_rvfi_mem_data_in_762,
  input  [31:0] io_rvfi_mem_data_in_763,
  input  [31:0] io_rvfi_mem_data_in_764,
  input  [31:0] io_rvfi_mem_data_in_765,
  input  [31:0] io_rvfi_mem_data_in_766,
  input  [31:0] io_rvfi_mem_data_in_767,
  input  [31:0] io_rvfi_mem_data_in_768,
  input  [31:0] io_rvfi_mem_data_in_769,
  input  [31:0] io_rvfi_mem_data_in_770,
  input  [31:0] io_rvfi_mem_data_in_771,
  input  [31:0] io_rvfi_mem_data_in_772,
  input  [31:0] io_rvfi_mem_data_in_773,
  input  [31:0] io_rvfi_mem_data_in_774,
  input  [31:0] io_rvfi_mem_data_in_775,
  input  [31:0] io_rvfi_mem_data_in_776,
  input  [31:0] io_rvfi_mem_data_in_777,
  input  [31:0] io_rvfi_mem_data_in_778,
  input  [31:0] io_rvfi_mem_data_in_779,
  input  [31:0] io_rvfi_mem_data_in_780,
  input  [31:0] io_rvfi_mem_data_in_781,
  input  [31:0] io_rvfi_mem_data_in_782,
  input  [31:0] io_rvfi_mem_data_in_783,
  input  [31:0] io_rvfi_mem_data_in_784,
  input  [31:0] io_rvfi_mem_data_in_785,
  input  [31:0] io_rvfi_mem_data_in_786,
  input  [31:0] io_rvfi_mem_data_in_787,
  input  [31:0] io_rvfi_mem_data_in_788,
  input  [31:0] io_rvfi_mem_data_in_789,
  input  [31:0] io_rvfi_mem_data_in_790,
  input  [31:0] io_rvfi_mem_data_in_791,
  input  [31:0] io_rvfi_mem_data_in_792,
  input  [31:0] io_rvfi_mem_data_in_793,
  input  [31:0] io_rvfi_mem_data_in_794,
  input  [31:0] io_rvfi_mem_data_in_795,
  input  [31:0] io_rvfi_mem_data_in_796,
  input  [31:0] io_rvfi_mem_data_in_797,
  input  [31:0] io_rvfi_mem_data_in_798,
  input  [31:0] io_rvfi_mem_data_in_799,
  input  [31:0] io_rvfi_mem_data_in_800,
  input  [31:0] io_rvfi_mem_data_in_801,
  input  [31:0] io_rvfi_mem_data_in_802,
  input  [31:0] io_rvfi_mem_data_in_803,
  input  [31:0] io_rvfi_mem_data_in_804,
  input  [31:0] io_rvfi_mem_data_in_805,
  input  [31:0] io_rvfi_mem_data_in_806,
  input  [31:0] io_rvfi_mem_data_in_807,
  input  [31:0] io_rvfi_mem_data_in_808,
  input  [31:0] io_rvfi_mem_data_in_809,
  input  [31:0] io_rvfi_mem_data_in_810,
  input  [31:0] io_rvfi_mem_data_in_811,
  input  [31:0] io_rvfi_mem_data_in_812,
  input  [31:0] io_rvfi_mem_data_in_813,
  input  [31:0] io_rvfi_mem_data_in_814,
  input  [31:0] io_rvfi_mem_data_in_815,
  input  [31:0] io_rvfi_mem_data_in_816,
  input  [31:0] io_rvfi_mem_data_in_817,
  input  [31:0] io_rvfi_mem_data_in_818,
  input  [31:0] io_rvfi_mem_data_in_819,
  input  [31:0] io_rvfi_mem_data_in_820,
  input  [31:0] io_rvfi_mem_data_in_821,
  input  [31:0] io_rvfi_mem_data_in_822,
  input  [31:0] io_rvfi_mem_data_in_823,
  input  [31:0] io_rvfi_mem_data_in_824,
  input  [31:0] io_rvfi_mem_data_in_825,
  input  [31:0] io_rvfi_mem_data_in_826,
  input  [31:0] io_rvfi_mem_data_in_827,
  input  [31:0] io_rvfi_mem_data_in_828,
  input  [31:0] io_rvfi_mem_data_in_829,
  input  [31:0] io_rvfi_mem_data_in_830,
  input  [31:0] io_rvfi_mem_data_in_831,
  input  [31:0] io_rvfi_mem_data_in_832,
  input  [31:0] io_rvfi_mem_data_in_833,
  input  [31:0] io_rvfi_mem_data_in_834,
  input  [31:0] io_rvfi_mem_data_in_835,
  input  [31:0] io_rvfi_mem_data_in_836,
  input  [31:0] io_rvfi_mem_data_in_837,
  input  [31:0] io_rvfi_mem_data_in_838,
  input  [31:0] io_rvfi_mem_data_in_839,
  input  [31:0] io_rvfi_mem_data_in_840,
  input  [31:0] io_rvfi_mem_data_in_841,
  input  [31:0] io_rvfi_mem_data_in_842,
  input  [31:0] io_rvfi_mem_data_in_843,
  input  [31:0] io_rvfi_mem_data_in_844,
  input  [31:0] io_rvfi_mem_data_in_845,
  input  [31:0] io_rvfi_mem_data_in_846,
  input  [31:0] io_rvfi_mem_data_in_847,
  input  [31:0] io_rvfi_mem_data_in_848,
  input  [31:0] io_rvfi_mem_data_in_849,
  input  [31:0] io_rvfi_mem_data_in_850,
  input  [31:0] io_rvfi_mem_data_in_851,
  input  [31:0] io_rvfi_mem_data_in_852,
  input  [31:0] io_rvfi_mem_data_in_853,
  input  [31:0] io_rvfi_mem_data_in_854,
  input  [31:0] io_rvfi_mem_data_in_855,
  input  [31:0] io_rvfi_mem_data_in_856,
  input  [31:0] io_rvfi_mem_data_in_857,
  input  [31:0] io_rvfi_mem_data_in_858,
  input  [31:0] io_rvfi_mem_data_in_859,
  input  [31:0] io_rvfi_mem_data_in_860,
  input  [31:0] io_rvfi_mem_data_in_861,
  input  [31:0] io_rvfi_mem_data_in_862,
  input  [31:0] io_rvfi_mem_data_in_863,
  input  [31:0] io_rvfi_mem_data_in_864,
  input  [31:0] io_rvfi_mem_data_in_865,
  input  [31:0] io_rvfi_mem_data_in_866,
  input  [31:0] io_rvfi_mem_data_in_867,
  input  [31:0] io_rvfi_mem_data_in_868,
  input  [31:0] io_rvfi_mem_data_in_869,
  input  [31:0] io_rvfi_mem_data_in_870,
  input  [31:0] io_rvfi_mem_data_in_871,
  input  [31:0] io_rvfi_mem_data_in_872,
  input  [31:0] io_rvfi_mem_data_in_873,
  input  [31:0] io_rvfi_mem_data_in_874,
  input  [31:0] io_rvfi_mem_data_in_875,
  input  [31:0] io_rvfi_mem_data_in_876,
  input  [31:0] io_rvfi_mem_data_in_877,
  input  [31:0] io_rvfi_mem_data_in_878,
  input  [31:0] io_rvfi_mem_data_in_879,
  input  [31:0] io_rvfi_mem_data_in_880,
  input  [31:0] io_rvfi_mem_data_in_881,
  input  [31:0] io_rvfi_mem_data_in_882,
  input  [31:0] io_rvfi_mem_data_in_883,
  input  [31:0] io_rvfi_mem_data_in_884,
  input  [31:0] io_rvfi_mem_data_in_885,
  input  [31:0] io_rvfi_mem_data_in_886,
  input  [31:0] io_rvfi_mem_data_in_887,
  input  [31:0] io_rvfi_mem_data_in_888,
  input  [31:0] io_rvfi_mem_data_in_889,
  input  [31:0] io_rvfi_mem_data_in_890,
  input  [31:0] io_rvfi_mem_data_in_891,
  input  [31:0] io_rvfi_mem_data_in_892,
  input  [31:0] io_rvfi_mem_data_in_893,
  input  [31:0] io_rvfi_mem_data_in_894,
  input  [31:0] io_rvfi_mem_data_in_895,
  input  [31:0] io_rvfi_mem_data_in_896,
  input  [31:0] io_rvfi_mem_data_in_897,
  input  [31:0] io_rvfi_mem_data_in_898,
  input  [31:0] io_rvfi_mem_data_in_899,
  input  [31:0] io_rvfi_mem_data_in_900,
  input  [31:0] io_rvfi_mem_data_in_901,
  input  [31:0] io_rvfi_mem_data_in_902,
  input  [31:0] io_rvfi_mem_data_in_903,
  input  [31:0] io_rvfi_mem_data_in_904,
  input  [31:0] io_rvfi_mem_data_in_905,
  input  [31:0] io_rvfi_mem_data_in_906,
  input  [31:0] io_rvfi_mem_data_in_907,
  input  [31:0] io_rvfi_mem_data_in_908,
  input  [31:0] io_rvfi_mem_data_in_909,
  input  [31:0] io_rvfi_mem_data_in_910,
  input  [31:0] io_rvfi_mem_data_in_911,
  input  [31:0] io_rvfi_mem_data_in_912,
  input  [31:0] io_rvfi_mem_data_in_913,
  input  [31:0] io_rvfi_mem_data_in_914,
  input  [31:0] io_rvfi_mem_data_in_915,
  input  [31:0] io_rvfi_mem_data_in_916,
  input  [31:0] io_rvfi_mem_data_in_917,
  input  [31:0] io_rvfi_mem_data_in_918,
  input  [31:0] io_rvfi_mem_data_in_919,
  input  [31:0] io_rvfi_mem_data_in_920,
  input  [31:0] io_rvfi_mem_data_in_921,
  input  [31:0] io_rvfi_mem_data_in_922,
  input  [31:0] io_rvfi_mem_data_in_923,
  input  [31:0] io_rvfi_mem_data_in_924,
  input  [31:0] io_rvfi_mem_data_in_925,
  input  [31:0] io_rvfi_mem_data_in_926,
  input  [31:0] io_rvfi_mem_data_in_927,
  input  [31:0] io_rvfi_mem_data_in_928,
  input  [31:0] io_rvfi_mem_data_in_929,
  input  [31:0] io_rvfi_mem_data_in_930,
  input  [31:0] io_rvfi_mem_data_in_931,
  input  [31:0] io_rvfi_mem_data_in_932,
  input  [31:0] io_rvfi_mem_data_in_933,
  input  [31:0] io_rvfi_mem_data_in_934,
  input  [31:0] io_rvfi_mem_data_in_935,
  input  [31:0] io_rvfi_mem_data_in_936,
  input  [31:0] io_rvfi_mem_data_in_937,
  input  [31:0] io_rvfi_mem_data_in_938,
  input  [31:0] io_rvfi_mem_data_in_939,
  input  [31:0] io_rvfi_mem_data_in_940,
  input  [31:0] io_rvfi_mem_data_in_941,
  input  [31:0] io_rvfi_mem_data_in_942,
  input  [31:0] io_rvfi_mem_data_in_943,
  input  [31:0] io_rvfi_mem_data_in_944,
  input  [31:0] io_rvfi_mem_data_in_945,
  input  [31:0] io_rvfi_mem_data_in_946,
  input  [31:0] io_rvfi_mem_data_in_947,
  input  [31:0] io_rvfi_mem_data_in_948,
  input  [31:0] io_rvfi_mem_data_in_949,
  input  [31:0] io_rvfi_mem_data_in_950,
  input  [31:0] io_rvfi_mem_data_in_951,
  input  [31:0] io_rvfi_mem_data_in_952,
  input  [31:0] io_rvfi_mem_data_in_953,
  input  [31:0] io_rvfi_mem_data_in_954,
  input  [31:0] io_rvfi_mem_data_in_955,
  input  [31:0] io_rvfi_mem_data_in_956,
  input  [31:0] io_rvfi_mem_data_in_957,
  input  [31:0] io_rvfi_mem_data_in_958,
  input  [31:0] io_rvfi_mem_data_in_959,
  input  [31:0] io_rvfi_mem_data_in_960,
  input  [31:0] io_rvfi_mem_data_in_961,
  input  [31:0] io_rvfi_mem_data_in_962,
  input  [31:0] io_rvfi_mem_data_in_963,
  input  [31:0] io_rvfi_mem_data_in_964,
  input  [31:0] io_rvfi_mem_data_in_965,
  input  [31:0] io_rvfi_mem_data_in_966,
  input  [31:0] io_rvfi_mem_data_in_967,
  input  [31:0] io_rvfi_mem_data_in_968,
  input  [31:0] io_rvfi_mem_data_in_969,
  input  [31:0] io_rvfi_mem_data_in_970,
  input  [31:0] io_rvfi_mem_data_in_971,
  input  [31:0] io_rvfi_mem_data_in_972,
  input  [31:0] io_rvfi_mem_data_in_973,
  input  [31:0] io_rvfi_mem_data_in_974,
  input  [31:0] io_rvfi_mem_data_in_975,
  input  [31:0] io_rvfi_mem_data_in_976,
  input  [31:0] io_rvfi_mem_data_in_977,
  input  [31:0] io_rvfi_mem_data_in_978,
  input  [31:0] io_rvfi_mem_data_in_979,
  input  [31:0] io_rvfi_mem_data_in_980,
  input  [31:0] io_rvfi_mem_data_in_981,
  input  [31:0] io_rvfi_mem_data_in_982,
  input  [31:0] io_rvfi_mem_data_in_983,
  input  [31:0] io_rvfi_mem_data_in_984,
  input  [31:0] io_rvfi_mem_data_in_985,
  input  [31:0] io_rvfi_mem_data_in_986,
  input  [31:0] io_rvfi_mem_data_in_987,
  input  [31:0] io_rvfi_mem_data_in_988,
  input  [31:0] io_rvfi_mem_data_in_989,
  input  [31:0] io_rvfi_mem_data_in_990,
  input  [31:0] io_rvfi_mem_data_in_991,
  input  [31:0] io_rvfi_mem_data_in_992,
  input  [31:0] io_rvfi_mem_data_in_993,
  input  [31:0] io_rvfi_mem_data_in_994,
  input  [31:0] io_rvfi_mem_data_in_995,
  input  [31:0] io_rvfi_mem_data_in_996,
  input  [31:0] io_rvfi_mem_data_in_997,
  input  [31:0] io_rvfi_mem_data_in_998,
  input  [31:0] io_rvfi_mem_data_in_999,
  input  [31:0] io_rvfi_mem_data_in_1000,
  input  [31:0] io_rvfi_mem_data_in_1001,
  input  [31:0] io_rvfi_mem_data_in_1002,
  input  [31:0] io_rvfi_mem_data_in_1003,
  input  [31:0] io_rvfi_mem_data_in_1004,
  input  [31:0] io_rvfi_mem_data_in_1005,
  input  [31:0] io_rvfi_mem_data_in_1006,
  input  [31:0] io_rvfi_mem_data_in_1007,
  input  [31:0] io_rvfi_mem_data_in_1008,
  input  [31:0] io_rvfi_mem_data_in_1009,
  input  [31:0] io_rvfi_mem_data_in_1010,
  input  [31:0] io_rvfi_mem_data_in_1011,
  input  [31:0] io_rvfi_mem_data_in_1012,
  input  [31:0] io_rvfi_mem_data_in_1013,
  input  [31:0] io_rvfi_mem_data_in_1014,
  input  [31:0] io_rvfi_mem_data_in_1015,
  input  [31:0] io_rvfi_mem_data_in_1016,
  input  [31:0] io_rvfi_mem_data_in_1017,
  input  [31:0] io_rvfi_mem_data_in_1018,
  input  [31:0] io_rvfi_mem_data_in_1019,
  input  [31:0] io_rvfi_mem_data_in_1020,
  input  [31:0] io_rvfi_mem_data_in_1021,
  input  [31:0] io_rvfi_mem_data_in_1022,
  input  [31:0] io_rvfi_mem_data_in_1023,
  output        io_rvfi_valid,
  output [31:0] io_rvfi_insn,
  output [63:0] io_rvfi_pc_rdata,
  output [63:0] io_rvfi_pc_wdata,
  output [4:0]  io_rvfi_rs1_addr,
  output [4:0]  io_rvfi_rs2_addr,
  output [63:0] io_rvfi_rs1_rdata,
  output [63:0] io_rvfi_rs2_rdata,
  output [4:0]  io_rvfi_rd_addr,
  output [63:0] io_rvfi_rd_wdata,
  output [31:0] io_rvfi_mem_addr,
  output [63:0] io_rvfi_mem_rdata,
  output [63:0] io_rvfi_mem_wdata,
  output [63:0] io_rvfi_regs_0,
  output [63:0] io_rvfi_regs_1,
  output [63:0] io_rvfi_regs_2,
  output [63:0] io_rvfi_regs_3,
  output [63:0] io_rvfi_regs_4,
  output [63:0] io_rvfi_regs_5,
  output [63:0] io_rvfi_regs_6,
  output [63:0] io_rvfi_regs_7,
  output [63:0] io_rvfi_regs_8,
  output [63:0] io_rvfi_regs_9,
  output [63:0] io_rvfi_regs_10,
  output [63:0] io_rvfi_regs_11,
  output [63:0] io_rvfi_regs_12,
  output [63:0] io_rvfi_regs_13,
  output [63:0] io_rvfi_regs_14,
  output [63:0] io_rvfi_regs_15,
  output [63:0] io_rvfi_regs_16,
  output [63:0] io_rvfi_regs_17,
  output [63:0] io_rvfi_regs_18,
  output [63:0] io_rvfi_regs_19,
  output [63:0] io_rvfi_regs_20,
  output [63:0] io_rvfi_regs_21,
  output [63:0] io_rvfi_regs_22,
  output [63:0] io_rvfi_regs_23,
  output [63:0] io_rvfi_regs_24,
  output [63:0] io_rvfi_regs_25,
  output [63:0] io_rvfi_regs_26,
  output [63:0] io_rvfi_regs_27,
  output [63:0] io_rvfi_regs_28,
  output [63:0] io_rvfi_regs_29,
  output [63:0] io_rvfi_regs_30,
  output [63:0] io_rvfi_regs_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [63:0] _RAND_1074;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] PC; // @[cpu.scala 42:19]
  reg [63:0] Regs_0; // @[cpu.scala 43:17]
  reg [63:0] Regs_1; // @[cpu.scala 43:17]
  reg [63:0] Regs_2; // @[cpu.scala 43:17]
  reg [63:0] Regs_3; // @[cpu.scala 43:17]
  reg [63:0] Regs_4; // @[cpu.scala 43:17]
  reg [63:0] Regs_5; // @[cpu.scala 43:17]
  reg [63:0] Regs_6; // @[cpu.scala 43:17]
  reg [63:0] Regs_7; // @[cpu.scala 43:17]
  reg [63:0] Regs_8; // @[cpu.scala 43:17]
  reg [63:0] Regs_9; // @[cpu.scala 43:17]
  reg [63:0] Regs_10; // @[cpu.scala 43:17]
  reg [63:0] Regs_11; // @[cpu.scala 43:17]
  reg [63:0] Regs_12; // @[cpu.scala 43:17]
  reg [63:0] Regs_13; // @[cpu.scala 43:17]
  reg [63:0] Regs_14; // @[cpu.scala 43:17]
  reg [63:0] Regs_15; // @[cpu.scala 43:17]
  reg [63:0] Regs_16; // @[cpu.scala 43:17]
  reg [63:0] Regs_17; // @[cpu.scala 43:17]
  reg [63:0] Regs_18; // @[cpu.scala 43:17]
  reg [63:0] Regs_19; // @[cpu.scala 43:17]
  reg [63:0] Regs_20; // @[cpu.scala 43:17]
  reg [63:0] Regs_21; // @[cpu.scala 43:17]
  reg [63:0] Regs_22; // @[cpu.scala 43:17]
  reg [63:0] Regs_23; // @[cpu.scala 43:17]
  reg [63:0] Regs_24; // @[cpu.scala 43:17]
  reg [63:0] Regs_25; // @[cpu.scala 43:17]
  reg [63:0] Regs_26; // @[cpu.scala 43:17]
  reg [63:0] Regs_27; // @[cpu.scala 43:17]
  reg [63:0] Regs_28; // @[cpu.scala 43:17]
  reg [63:0] Regs_29; // @[cpu.scala 43:17]
  reg [63:0] Regs_30; // @[cpu.scala 43:17]
  reg [63:0] Regs_31; // @[cpu.scala 43:17]
  reg [63:0] IDEXA; // @[cpu.scala 44:58]
  reg [63:0] IDEXB; // @[cpu.scala 44:58]
  reg [63:0] EXMEMB; // @[cpu.scala 44:58]
  reg [63:0] EXMEMALUOut; // @[cpu.scala 44:58]
  reg [63:0] MEMWBValue; // @[cpu.scala 44:58]
  reg [31:0] DMemory_0; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1; // @[cpu.scala 46:20]
  reg [31:0] DMemory_2; // @[cpu.scala 46:20]
  reg [31:0] DMemory_3; // @[cpu.scala 46:20]
  reg [31:0] DMemory_4; // @[cpu.scala 46:20]
  reg [31:0] DMemory_5; // @[cpu.scala 46:20]
  reg [31:0] DMemory_6; // @[cpu.scala 46:20]
  reg [31:0] DMemory_7; // @[cpu.scala 46:20]
  reg [31:0] DMemory_8; // @[cpu.scala 46:20]
  reg [31:0] DMemory_9; // @[cpu.scala 46:20]
  reg [31:0] DMemory_10; // @[cpu.scala 46:20]
  reg [31:0] DMemory_11; // @[cpu.scala 46:20]
  reg [31:0] DMemory_12; // @[cpu.scala 46:20]
  reg [31:0] DMemory_13; // @[cpu.scala 46:20]
  reg [31:0] DMemory_14; // @[cpu.scala 46:20]
  reg [31:0] DMemory_15; // @[cpu.scala 46:20]
  reg [31:0] DMemory_16; // @[cpu.scala 46:20]
  reg [31:0] DMemory_17; // @[cpu.scala 46:20]
  reg [31:0] DMemory_18; // @[cpu.scala 46:20]
  reg [31:0] DMemory_19; // @[cpu.scala 46:20]
  reg [31:0] DMemory_20; // @[cpu.scala 46:20]
  reg [31:0] DMemory_21; // @[cpu.scala 46:20]
  reg [31:0] DMemory_22; // @[cpu.scala 46:20]
  reg [31:0] DMemory_23; // @[cpu.scala 46:20]
  reg [31:0] DMemory_24; // @[cpu.scala 46:20]
  reg [31:0] DMemory_25; // @[cpu.scala 46:20]
  reg [31:0] DMemory_26; // @[cpu.scala 46:20]
  reg [31:0] DMemory_27; // @[cpu.scala 46:20]
  reg [31:0] DMemory_28; // @[cpu.scala 46:20]
  reg [31:0] DMemory_29; // @[cpu.scala 46:20]
  reg [31:0] DMemory_30; // @[cpu.scala 46:20]
  reg [31:0] DMemory_31; // @[cpu.scala 46:20]
  reg [31:0] DMemory_32; // @[cpu.scala 46:20]
  reg [31:0] DMemory_33; // @[cpu.scala 46:20]
  reg [31:0] DMemory_34; // @[cpu.scala 46:20]
  reg [31:0] DMemory_35; // @[cpu.scala 46:20]
  reg [31:0] DMemory_36; // @[cpu.scala 46:20]
  reg [31:0] DMemory_37; // @[cpu.scala 46:20]
  reg [31:0] DMemory_38; // @[cpu.scala 46:20]
  reg [31:0] DMemory_39; // @[cpu.scala 46:20]
  reg [31:0] DMemory_40; // @[cpu.scala 46:20]
  reg [31:0] DMemory_41; // @[cpu.scala 46:20]
  reg [31:0] DMemory_42; // @[cpu.scala 46:20]
  reg [31:0] DMemory_43; // @[cpu.scala 46:20]
  reg [31:0] DMemory_44; // @[cpu.scala 46:20]
  reg [31:0] DMemory_45; // @[cpu.scala 46:20]
  reg [31:0] DMemory_46; // @[cpu.scala 46:20]
  reg [31:0] DMemory_47; // @[cpu.scala 46:20]
  reg [31:0] DMemory_48; // @[cpu.scala 46:20]
  reg [31:0] DMemory_49; // @[cpu.scala 46:20]
  reg [31:0] DMemory_50; // @[cpu.scala 46:20]
  reg [31:0] DMemory_51; // @[cpu.scala 46:20]
  reg [31:0] DMemory_52; // @[cpu.scala 46:20]
  reg [31:0] DMemory_53; // @[cpu.scala 46:20]
  reg [31:0] DMemory_54; // @[cpu.scala 46:20]
  reg [31:0] DMemory_55; // @[cpu.scala 46:20]
  reg [31:0] DMemory_56; // @[cpu.scala 46:20]
  reg [31:0] DMemory_57; // @[cpu.scala 46:20]
  reg [31:0] DMemory_58; // @[cpu.scala 46:20]
  reg [31:0] DMemory_59; // @[cpu.scala 46:20]
  reg [31:0] DMemory_60; // @[cpu.scala 46:20]
  reg [31:0] DMemory_61; // @[cpu.scala 46:20]
  reg [31:0] DMemory_62; // @[cpu.scala 46:20]
  reg [31:0] DMemory_63; // @[cpu.scala 46:20]
  reg [31:0] DMemory_64; // @[cpu.scala 46:20]
  reg [31:0] DMemory_65; // @[cpu.scala 46:20]
  reg [31:0] DMemory_66; // @[cpu.scala 46:20]
  reg [31:0] DMemory_67; // @[cpu.scala 46:20]
  reg [31:0] DMemory_68; // @[cpu.scala 46:20]
  reg [31:0] DMemory_69; // @[cpu.scala 46:20]
  reg [31:0] DMemory_70; // @[cpu.scala 46:20]
  reg [31:0] DMemory_71; // @[cpu.scala 46:20]
  reg [31:0] DMemory_72; // @[cpu.scala 46:20]
  reg [31:0] DMemory_73; // @[cpu.scala 46:20]
  reg [31:0] DMemory_74; // @[cpu.scala 46:20]
  reg [31:0] DMemory_75; // @[cpu.scala 46:20]
  reg [31:0] DMemory_76; // @[cpu.scala 46:20]
  reg [31:0] DMemory_77; // @[cpu.scala 46:20]
  reg [31:0] DMemory_78; // @[cpu.scala 46:20]
  reg [31:0] DMemory_79; // @[cpu.scala 46:20]
  reg [31:0] DMemory_80; // @[cpu.scala 46:20]
  reg [31:0] DMemory_81; // @[cpu.scala 46:20]
  reg [31:0] DMemory_82; // @[cpu.scala 46:20]
  reg [31:0] DMemory_83; // @[cpu.scala 46:20]
  reg [31:0] DMemory_84; // @[cpu.scala 46:20]
  reg [31:0] DMemory_85; // @[cpu.scala 46:20]
  reg [31:0] DMemory_86; // @[cpu.scala 46:20]
  reg [31:0] DMemory_87; // @[cpu.scala 46:20]
  reg [31:0] DMemory_88; // @[cpu.scala 46:20]
  reg [31:0] DMemory_89; // @[cpu.scala 46:20]
  reg [31:0] DMemory_90; // @[cpu.scala 46:20]
  reg [31:0] DMemory_91; // @[cpu.scala 46:20]
  reg [31:0] DMemory_92; // @[cpu.scala 46:20]
  reg [31:0] DMemory_93; // @[cpu.scala 46:20]
  reg [31:0] DMemory_94; // @[cpu.scala 46:20]
  reg [31:0] DMemory_95; // @[cpu.scala 46:20]
  reg [31:0] DMemory_96; // @[cpu.scala 46:20]
  reg [31:0] DMemory_97; // @[cpu.scala 46:20]
  reg [31:0] DMemory_98; // @[cpu.scala 46:20]
  reg [31:0] DMemory_99; // @[cpu.scala 46:20]
  reg [31:0] DMemory_100; // @[cpu.scala 46:20]
  reg [31:0] DMemory_101; // @[cpu.scala 46:20]
  reg [31:0] DMemory_102; // @[cpu.scala 46:20]
  reg [31:0] DMemory_103; // @[cpu.scala 46:20]
  reg [31:0] DMemory_104; // @[cpu.scala 46:20]
  reg [31:0] DMemory_105; // @[cpu.scala 46:20]
  reg [31:0] DMemory_106; // @[cpu.scala 46:20]
  reg [31:0] DMemory_107; // @[cpu.scala 46:20]
  reg [31:0] DMemory_108; // @[cpu.scala 46:20]
  reg [31:0] DMemory_109; // @[cpu.scala 46:20]
  reg [31:0] DMemory_110; // @[cpu.scala 46:20]
  reg [31:0] DMemory_111; // @[cpu.scala 46:20]
  reg [31:0] DMemory_112; // @[cpu.scala 46:20]
  reg [31:0] DMemory_113; // @[cpu.scala 46:20]
  reg [31:0] DMemory_114; // @[cpu.scala 46:20]
  reg [31:0] DMemory_115; // @[cpu.scala 46:20]
  reg [31:0] DMemory_116; // @[cpu.scala 46:20]
  reg [31:0] DMemory_117; // @[cpu.scala 46:20]
  reg [31:0] DMemory_118; // @[cpu.scala 46:20]
  reg [31:0] DMemory_119; // @[cpu.scala 46:20]
  reg [31:0] DMemory_120; // @[cpu.scala 46:20]
  reg [31:0] DMemory_121; // @[cpu.scala 46:20]
  reg [31:0] DMemory_122; // @[cpu.scala 46:20]
  reg [31:0] DMemory_123; // @[cpu.scala 46:20]
  reg [31:0] DMemory_124; // @[cpu.scala 46:20]
  reg [31:0] DMemory_125; // @[cpu.scala 46:20]
  reg [31:0] DMemory_126; // @[cpu.scala 46:20]
  reg [31:0] DMemory_127; // @[cpu.scala 46:20]
  reg [31:0] DMemory_128; // @[cpu.scala 46:20]
  reg [31:0] DMemory_129; // @[cpu.scala 46:20]
  reg [31:0] DMemory_130; // @[cpu.scala 46:20]
  reg [31:0] DMemory_131; // @[cpu.scala 46:20]
  reg [31:0] DMemory_132; // @[cpu.scala 46:20]
  reg [31:0] DMemory_133; // @[cpu.scala 46:20]
  reg [31:0] DMemory_134; // @[cpu.scala 46:20]
  reg [31:0] DMemory_135; // @[cpu.scala 46:20]
  reg [31:0] DMemory_136; // @[cpu.scala 46:20]
  reg [31:0] DMemory_137; // @[cpu.scala 46:20]
  reg [31:0] DMemory_138; // @[cpu.scala 46:20]
  reg [31:0] DMemory_139; // @[cpu.scala 46:20]
  reg [31:0] DMemory_140; // @[cpu.scala 46:20]
  reg [31:0] DMemory_141; // @[cpu.scala 46:20]
  reg [31:0] DMemory_142; // @[cpu.scala 46:20]
  reg [31:0] DMemory_143; // @[cpu.scala 46:20]
  reg [31:0] DMemory_144; // @[cpu.scala 46:20]
  reg [31:0] DMemory_145; // @[cpu.scala 46:20]
  reg [31:0] DMemory_146; // @[cpu.scala 46:20]
  reg [31:0] DMemory_147; // @[cpu.scala 46:20]
  reg [31:0] DMemory_148; // @[cpu.scala 46:20]
  reg [31:0] DMemory_149; // @[cpu.scala 46:20]
  reg [31:0] DMemory_150; // @[cpu.scala 46:20]
  reg [31:0] DMemory_151; // @[cpu.scala 46:20]
  reg [31:0] DMemory_152; // @[cpu.scala 46:20]
  reg [31:0] DMemory_153; // @[cpu.scala 46:20]
  reg [31:0] DMemory_154; // @[cpu.scala 46:20]
  reg [31:0] DMemory_155; // @[cpu.scala 46:20]
  reg [31:0] DMemory_156; // @[cpu.scala 46:20]
  reg [31:0] DMemory_157; // @[cpu.scala 46:20]
  reg [31:0] DMemory_158; // @[cpu.scala 46:20]
  reg [31:0] DMemory_159; // @[cpu.scala 46:20]
  reg [31:0] DMemory_160; // @[cpu.scala 46:20]
  reg [31:0] DMemory_161; // @[cpu.scala 46:20]
  reg [31:0] DMemory_162; // @[cpu.scala 46:20]
  reg [31:0] DMemory_163; // @[cpu.scala 46:20]
  reg [31:0] DMemory_164; // @[cpu.scala 46:20]
  reg [31:0] DMemory_165; // @[cpu.scala 46:20]
  reg [31:0] DMemory_166; // @[cpu.scala 46:20]
  reg [31:0] DMemory_167; // @[cpu.scala 46:20]
  reg [31:0] DMemory_168; // @[cpu.scala 46:20]
  reg [31:0] DMemory_169; // @[cpu.scala 46:20]
  reg [31:0] DMemory_170; // @[cpu.scala 46:20]
  reg [31:0] DMemory_171; // @[cpu.scala 46:20]
  reg [31:0] DMemory_172; // @[cpu.scala 46:20]
  reg [31:0] DMemory_173; // @[cpu.scala 46:20]
  reg [31:0] DMemory_174; // @[cpu.scala 46:20]
  reg [31:0] DMemory_175; // @[cpu.scala 46:20]
  reg [31:0] DMemory_176; // @[cpu.scala 46:20]
  reg [31:0] DMemory_177; // @[cpu.scala 46:20]
  reg [31:0] DMemory_178; // @[cpu.scala 46:20]
  reg [31:0] DMemory_179; // @[cpu.scala 46:20]
  reg [31:0] DMemory_180; // @[cpu.scala 46:20]
  reg [31:0] DMemory_181; // @[cpu.scala 46:20]
  reg [31:0] DMemory_182; // @[cpu.scala 46:20]
  reg [31:0] DMemory_183; // @[cpu.scala 46:20]
  reg [31:0] DMemory_184; // @[cpu.scala 46:20]
  reg [31:0] DMemory_185; // @[cpu.scala 46:20]
  reg [31:0] DMemory_186; // @[cpu.scala 46:20]
  reg [31:0] DMemory_187; // @[cpu.scala 46:20]
  reg [31:0] DMemory_188; // @[cpu.scala 46:20]
  reg [31:0] DMemory_189; // @[cpu.scala 46:20]
  reg [31:0] DMemory_190; // @[cpu.scala 46:20]
  reg [31:0] DMemory_191; // @[cpu.scala 46:20]
  reg [31:0] DMemory_192; // @[cpu.scala 46:20]
  reg [31:0] DMemory_193; // @[cpu.scala 46:20]
  reg [31:0] DMemory_194; // @[cpu.scala 46:20]
  reg [31:0] DMemory_195; // @[cpu.scala 46:20]
  reg [31:0] DMemory_196; // @[cpu.scala 46:20]
  reg [31:0] DMemory_197; // @[cpu.scala 46:20]
  reg [31:0] DMemory_198; // @[cpu.scala 46:20]
  reg [31:0] DMemory_199; // @[cpu.scala 46:20]
  reg [31:0] DMemory_200; // @[cpu.scala 46:20]
  reg [31:0] DMemory_201; // @[cpu.scala 46:20]
  reg [31:0] DMemory_202; // @[cpu.scala 46:20]
  reg [31:0] DMemory_203; // @[cpu.scala 46:20]
  reg [31:0] DMemory_204; // @[cpu.scala 46:20]
  reg [31:0] DMemory_205; // @[cpu.scala 46:20]
  reg [31:0] DMemory_206; // @[cpu.scala 46:20]
  reg [31:0] DMemory_207; // @[cpu.scala 46:20]
  reg [31:0] DMemory_208; // @[cpu.scala 46:20]
  reg [31:0] DMemory_209; // @[cpu.scala 46:20]
  reg [31:0] DMemory_210; // @[cpu.scala 46:20]
  reg [31:0] DMemory_211; // @[cpu.scala 46:20]
  reg [31:0] DMemory_212; // @[cpu.scala 46:20]
  reg [31:0] DMemory_213; // @[cpu.scala 46:20]
  reg [31:0] DMemory_214; // @[cpu.scala 46:20]
  reg [31:0] DMemory_215; // @[cpu.scala 46:20]
  reg [31:0] DMemory_216; // @[cpu.scala 46:20]
  reg [31:0] DMemory_217; // @[cpu.scala 46:20]
  reg [31:0] DMemory_218; // @[cpu.scala 46:20]
  reg [31:0] DMemory_219; // @[cpu.scala 46:20]
  reg [31:0] DMemory_220; // @[cpu.scala 46:20]
  reg [31:0] DMemory_221; // @[cpu.scala 46:20]
  reg [31:0] DMemory_222; // @[cpu.scala 46:20]
  reg [31:0] DMemory_223; // @[cpu.scala 46:20]
  reg [31:0] DMemory_224; // @[cpu.scala 46:20]
  reg [31:0] DMemory_225; // @[cpu.scala 46:20]
  reg [31:0] DMemory_226; // @[cpu.scala 46:20]
  reg [31:0] DMemory_227; // @[cpu.scala 46:20]
  reg [31:0] DMemory_228; // @[cpu.scala 46:20]
  reg [31:0] DMemory_229; // @[cpu.scala 46:20]
  reg [31:0] DMemory_230; // @[cpu.scala 46:20]
  reg [31:0] DMemory_231; // @[cpu.scala 46:20]
  reg [31:0] DMemory_232; // @[cpu.scala 46:20]
  reg [31:0] DMemory_233; // @[cpu.scala 46:20]
  reg [31:0] DMemory_234; // @[cpu.scala 46:20]
  reg [31:0] DMemory_235; // @[cpu.scala 46:20]
  reg [31:0] DMemory_236; // @[cpu.scala 46:20]
  reg [31:0] DMemory_237; // @[cpu.scala 46:20]
  reg [31:0] DMemory_238; // @[cpu.scala 46:20]
  reg [31:0] DMemory_239; // @[cpu.scala 46:20]
  reg [31:0] DMemory_240; // @[cpu.scala 46:20]
  reg [31:0] DMemory_241; // @[cpu.scala 46:20]
  reg [31:0] DMemory_242; // @[cpu.scala 46:20]
  reg [31:0] DMemory_243; // @[cpu.scala 46:20]
  reg [31:0] DMemory_244; // @[cpu.scala 46:20]
  reg [31:0] DMemory_245; // @[cpu.scala 46:20]
  reg [31:0] DMemory_246; // @[cpu.scala 46:20]
  reg [31:0] DMemory_247; // @[cpu.scala 46:20]
  reg [31:0] DMemory_248; // @[cpu.scala 46:20]
  reg [31:0] DMemory_249; // @[cpu.scala 46:20]
  reg [31:0] DMemory_250; // @[cpu.scala 46:20]
  reg [31:0] DMemory_251; // @[cpu.scala 46:20]
  reg [31:0] DMemory_252; // @[cpu.scala 46:20]
  reg [31:0] DMemory_253; // @[cpu.scala 46:20]
  reg [31:0] DMemory_254; // @[cpu.scala 46:20]
  reg [31:0] DMemory_255; // @[cpu.scala 46:20]
  reg [31:0] DMemory_256; // @[cpu.scala 46:20]
  reg [31:0] DMemory_257; // @[cpu.scala 46:20]
  reg [31:0] DMemory_258; // @[cpu.scala 46:20]
  reg [31:0] DMemory_259; // @[cpu.scala 46:20]
  reg [31:0] DMemory_260; // @[cpu.scala 46:20]
  reg [31:0] DMemory_261; // @[cpu.scala 46:20]
  reg [31:0] DMemory_262; // @[cpu.scala 46:20]
  reg [31:0] DMemory_263; // @[cpu.scala 46:20]
  reg [31:0] DMemory_264; // @[cpu.scala 46:20]
  reg [31:0] DMemory_265; // @[cpu.scala 46:20]
  reg [31:0] DMemory_266; // @[cpu.scala 46:20]
  reg [31:0] DMemory_267; // @[cpu.scala 46:20]
  reg [31:0] DMemory_268; // @[cpu.scala 46:20]
  reg [31:0] DMemory_269; // @[cpu.scala 46:20]
  reg [31:0] DMemory_270; // @[cpu.scala 46:20]
  reg [31:0] DMemory_271; // @[cpu.scala 46:20]
  reg [31:0] DMemory_272; // @[cpu.scala 46:20]
  reg [31:0] DMemory_273; // @[cpu.scala 46:20]
  reg [31:0] DMemory_274; // @[cpu.scala 46:20]
  reg [31:0] DMemory_275; // @[cpu.scala 46:20]
  reg [31:0] DMemory_276; // @[cpu.scala 46:20]
  reg [31:0] DMemory_277; // @[cpu.scala 46:20]
  reg [31:0] DMemory_278; // @[cpu.scala 46:20]
  reg [31:0] DMemory_279; // @[cpu.scala 46:20]
  reg [31:0] DMemory_280; // @[cpu.scala 46:20]
  reg [31:0] DMemory_281; // @[cpu.scala 46:20]
  reg [31:0] DMemory_282; // @[cpu.scala 46:20]
  reg [31:0] DMemory_283; // @[cpu.scala 46:20]
  reg [31:0] DMemory_284; // @[cpu.scala 46:20]
  reg [31:0] DMemory_285; // @[cpu.scala 46:20]
  reg [31:0] DMemory_286; // @[cpu.scala 46:20]
  reg [31:0] DMemory_287; // @[cpu.scala 46:20]
  reg [31:0] DMemory_288; // @[cpu.scala 46:20]
  reg [31:0] DMemory_289; // @[cpu.scala 46:20]
  reg [31:0] DMemory_290; // @[cpu.scala 46:20]
  reg [31:0] DMemory_291; // @[cpu.scala 46:20]
  reg [31:0] DMemory_292; // @[cpu.scala 46:20]
  reg [31:0] DMemory_293; // @[cpu.scala 46:20]
  reg [31:0] DMemory_294; // @[cpu.scala 46:20]
  reg [31:0] DMemory_295; // @[cpu.scala 46:20]
  reg [31:0] DMemory_296; // @[cpu.scala 46:20]
  reg [31:0] DMemory_297; // @[cpu.scala 46:20]
  reg [31:0] DMemory_298; // @[cpu.scala 46:20]
  reg [31:0] DMemory_299; // @[cpu.scala 46:20]
  reg [31:0] DMemory_300; // @[cpu.scala 46:20]
  reg [31:0] DMemory_301; // @[cpu.scala 46:20]
  reg [31:0] DMemory_302; // @[cpu.scala 46:20]
  reg [31:0] DMemory_303; // @[cpu.scala 46:20]
  reg [31:0] DMemory_304; // @[cpu.scala 46:20]
  reg [31:0] DMemory_305; // @[cpu.scala 46:20]
  reg [31:0] DMemory_306; // @[cpu.scala 46:20]
  reg [31:0] DMemory_307; // @[cpu.scala 46:20]
  reg [31:0] DMemory_308; // @[cpu.scala 46:20]
  reg [31:0] DMemory_309; // @[cpu.scala 46:20]
  reg [31:0] DMemory_310; // @[cpu.scala 46:20]
  reg [31:0] DMemory_311; // @[cpu.scala 46:20]
  reg [31:0] DMemory_312; // @[cpu.scala 46:20]
  reg [31:0] DMemory_313; // @[cpu.scala 46:20]
  reg [31:0] DMemory_314; // @[cpu.scala 46:20]
  reg [31:0] DMemory_315; // @[cpu.scala 46:20]
  reg [31:0] DMemory_316; // @[cpu.scala 46:20]
  reg [31:0] DMemory_317; // @[cpu.scala 46:20]
  reg [31:0] DMemory_318; // @[cpu.scala 46:20]
  reg [31:0] DMemory_319; // @[cpu.scala 46:20]
  reg [31:0] DMemory_320; // @[cpu.scala 46:20]
  reg [31:0] DMemory_321; // @[cpu.scala 46:20]
  reg [31:0] DMemory_322; // @[cpu.scala 46:20]
  reg [31:0] DMemory_323; // @[cpu.scala 46:20]
  reg [31:0] DMemory_324; // @[cpu.scala 46:20]
  reg [31:0] DMemory_325; // @[cpu.scala 46:20]
  reg [31:0] DMemory_326; // @[cpu.scala 46:20]
  reg [31:0] DMemory_327; // @[cpu.scala 46:20]
  reg [31:0] DMemory_328; // @[cpu.scala 46:20]
  reg [31:0] DMemory_329; // @[cpu.scala 46:20]
  reg [31:0] DMemory_330; // @[cpu.scala 46:20]
  reg [31:0] DMemory_331; // @[cpu.scala 46:20]
  reg [31:0] DMemory_332; // @[cpu.scala 46:20]
  reg [31:0] DMemory_333; // @[cpu.scala 46:20]
  reg [31:0] DMemory_334; // @[cpu.scala 46:20]
  reg [31:0] DMemory_335; // @[cpu.scala 46:20]
  reg [31:0] DMemory_336; // @[cpu.scala 46:20]
  reg [31:0] DMemory_337; // @[cpu.scala 46:20]
  reg [31:0] DMemory_338; // @[cpu.scala 46:20]
  reg [31:0] DMemory_339; // @[cpu.scala 46:20]
  reg [31:0] DMemory_340; // @[cpu.scala 46:20]
  reg [31:0] DMemory_341; // @[cpu.scala 46:20]
  reg [31:0] DMemory_342; // @[cpu.scala 46:20]
  reg [31:0] DMemory_343; // @[cpu.scala 46:20]
  reg [31:0] DMemory_344; // @[cpu.scala 46:20]
  reg [31:0] DMemory_345; // @[cpu.scala 46:20]
  reg [31:0] DMemory_346; // @[cpu.scala 46:20]
  reg [31:0] DMemory_347; // @[cpu.scala 46:20]
  reg [31:0] DMemory_348; // @[cpu.scala 46:20]
  reg [31:0] DMemory_349; // @[cpu.scala 46:20]
  reg [31:0] DMemory_350; // @[cpu.scala 46:20]
  reg [31:0] DMemory_351; // @[cpu.scala 46:20]
  reg [31:0] DMemory_352; // @[cpu.scala 46:20]
  reg [31:0] DMemory_353; // @[cpu.scala 46:20]
  reg [31:0] DMemory_354; // @[cpu.scala 46:20]
  reg [31:0] DMemory_355; // @[cpu.scala 46:20]
  reg [31:0] DMemory_356; // @[cpu.scala 46:20]
  reg [31:0] DMemory_357; // @[cpu.scala 46:20]
  reg [31:0] DMemory_358; // @[cpu.scala 46:20]
  reg [31:0] DMemory_359; // @[cpu.scala 46:20]
  reg [31:0] DMemory_360; // @[cpu.scala 46:20]
  reg [31:0] DMemory_361; // @[cpu.scala 46:20]
  reg [31:0] DMemory_362; // @[cpu.scala 46:20]
  reg [31:0] DMemory_363; // @[cpu.scala 46:20]
  reg [31:0] DMemory_364; // @[cpu.scala 46:20]
  reg [31:0] DMemory_365; // @[cpu.scala 46:20]
  reg [31:0] DMemory_366; // @[cpu.scala 46:20]
  reg [31:0] DMemory_367; // @[cpu.scala 46:20]
  reg [31:0] DMemory_368; // @[cpu.scala 46:20]
  reg [31:0] DMemory_369; // @[cpu.scala 46:20]
  reg [31:0] DMemory_370; // @[cpu.scala 46:20]
  reg [31:0] DMemory_371; // @[cpu.scala 46:20]
  reg [31:0] DMemory_372; // @[cpu.scala 46:20]
  reg [31:0] DMemory_373; // @[cpu.scala 46:20]
  reg [31:0] DMemory_374; // @[cpu.scala 46:20]
  reg [31:0] DMemory_375; // @[cpu.scala 46:20]
  reg [31:0] DMemory_376; // @[cpu.scala 46:20]
  reg [31:0] DMemory_377; // @[cpu.scala 46:20]
  reg [31:0] DMemory_378; // @[cpu.scala 46:20]
  reg [31:0] DMemory_379; // @[cpu.scala 46:20]
  reg [31:0] DMemory_380; // @[cpu.scala 46:20]
  reg [31:0] DMemory_381; // @[cpu.scala 46:20]
  reg [31:0] DMemory_382; // @[cpu.scala 46:20]
  reg [31:0] DMemory_383; // @[cpu.scala 46:20]
  reg [31:0] DMemory_384; // @[cpu.scala 46:20]
  reg [31:0] DMemory_385; // @[cpu.scala 46:20]
  reg [31:0] DMemory_386; // @[cpu.scala 46:20]
  reg [31:0] DMemory_387; // @[cpu.scala 46:20]
  reg [31:0] DMemory_388; // @[cpu.scala 46:20]
  reg [31:0] DMemory_389; // @[cpu.scala 46:20]
  reg [31:0] DMemory_390; // @[cpu.scala 46:20]
  reg [31:0] DMemory_391; // @[cpu.scala 46:20]
  reg [31:0] DMemory_392; // @[cpu.scala 46:20]
  reg [31:0] DMemory_393; // @[cpu.scala 46:20]
  reg [31:0] DMemory_394; // @[cpu.scala 46:20]
  reg [31:0] DMemory_395; // @[cpu.scala 46:20]
  reg [31:0] DMemory_396; // @[cpu.scala 46:20]
  reg [31:0] DMemory_397; // @[cpu.scala 46:20]
  reg [31:0] DMemory_398; // @[cpu.scala 46:20]
  reg [31:0] DMemory_399; // @[cpu.scala 46:20]
  reg [31:0] DMemory_400; // @[cpu.scala 46:20]
  reg [31:0] DMemory_401; // @[cpu.scala 46:20]
  reg [31:0] DMemory_402; // @[cpu.scala 46:20]
  reg [31:0] DMemory_403; // @[cpu.scala 46:20]
  reg [31:0] DMemory_404; // @[cpu.scala 46:20]
  reg [31:0] DMemory_405; // @[cpu.scala 46:20]
  reg [31:0] DMemory_406; // @[cpu.scala 46:20]
  reg [31:0] DMemory_407; // @[cpu.scala 46:20]
  reg [31:0] DMemory_408; // @[cpu.scala 46:20]
  reg [31:0] DMemory_409; // @[cpu.scala 46:20]
  reg [31:0] DMemory_410; // @[cpu.scala 46:20]
  reg [31:0] DMemory_411; // @[cpu.scala 46:20]
  reg [31:0] DMemory_412; // @[cpu.scala 46:20]
  reg [31:0] DMemory_413; // @[cpu.scala 46:20]
  reg [31:0] DMemory_414; // @[cpu.scala 46:20]
  reg [31:0] DMemory_415; // @[cpu.scala 46:20]
  reg [31:0] DMemory_416; // @[cpu.scala 46:20]
  reg [31:0] DMemory_417; // @[cpu.scala 46:20]
  reg [31:0] DMemory_418; // @[cpu.scala 46:20]
  reg [31:0] DMemory_419; // @[cpu.scala 46:20]
  reg [31:0] DMemory_420; // @[cpu.scala 46:20]
  reg [31:0] DMemory_421; // @[cpu.scala 46:20]
  reg [31:0] DMemory_422; // @[cpu.scala 46:20]
  reg [31:0] DMemory_423; // @[cpu.scala 46:20]
  reg [31:0] DMemory_424; // @[cpu.scala 46:20]
  reg [31:0] DMemory_425; // @[cpu.scala 46:20]
  reg [31:0] DMemory_426; // @[cpu.scala 46:20]
  reg [31:0] DMemory_427; // @[cpu.scala 46:20]
  reg [31:0] DMemory_428; // @[cpu.scala 46:20]
  reg [31:0] DMemory_429; // @[cpu.scala 46:20]
  reg [31:0] DMemory_430; // @[cpu.scala 46:20]
  reg [31:0] DMemory_431; // @[cpu.scala 46:20]
  reg [31:0] DMemory_432; // @[cpu.scala 46:20]
  reg [31:0] DMemory_433; // @[cpu.scala 46:20]
  reg [31:0] DMemory_434; // @[cpu.scala 46:20]
  reg [31:0] DMemory_435; // @[cpu.scala 46:20]
  reg [31:0] DMemory_436; // @[cpu.scala 46:20]
  reg [31:0] DMemory_437; // @[cpu.scala 46:20]
  reg [31:0] DMemory_438; // @[cpu.scala 46:20]
  reg [31:0] DMemory_439; // @[cpu.scala 46:20]
  reg [31:0] DMemory_440; // @[cpu.scala 46:20]
  reg [31:0] DMemory_441; // @[cpu.scala 46:20]
  reg [31:0] DMemory_442; // @[cpu.scala 46:20]
  reg [31:0] DMemory_443; // @[cpu.scala 46:20]
  reg [31:0] DMemory_444; // @[cpu.scala 46:20]
  reg [31:0] DMemory_445; // @[cpu.scala 46:20]
  reg [31:0] DMemory_446; // @[cpu.scala 46:20]
  reg [31:0] DMemory_447; // @[cpu.scala 46:20]
  reg [31:0] DMemory_448; // @[cpu.scala 46:20]
  reg [31:0] DMemory_449; // @[cpu.scala 46:20]
  reg [31:0] DMemory_450; // @[cpu.scala 46:20]
  reg [31:0] DMemory_451; // @[cpu.scala 46:20]
  reg [31:0] DMemory_452; // @[cpu.scala 46:20]
  reg [31:0] DMemory_453; // @[cpu.scala 46:20]
  reg [31:0] DMemory_454; // @[cpu.scala 46:20]
  reg [31:0] DMemory_455; // @[cpu.scala 46:20]
  reg [31:0] DMemory_456; // @[cpu.scala 46:20]
  reg [31:0] DMemory_457; // @[cpu.scala 46:20]
  reg [31:0] DMemory_458; // @[cpu.scala 46:20]
  reg [31:0] DMemory_459; // @[cpu.scala 46:20]
  reg [31:0] DMemory_460; // @[cpu.scala 46:20]
  reg [31:0] DMemory_461; // @[cpu.scala 46:20]
  reg [31:0] DMemory_462; // @[cpu.scala 46:20]
  reg [31:0] DMemory_463; // @[cpu.scala 46:20]
  reg [31:0] DMemory_464; // @[cpu.scala 46:20]
  reg [31:0] DMemory_465; // @[cpu.scala 46:20]
  reg [31:0] DMemory_466; // @[cpu.scala 46:20]
  reg [31:0] DMemory_467; // @[cpu.scala 46:20]
  reg [31:0] DMemory_468; // @[cpu.scala 46:20]
  reg [31:0] DMemory_469; // @[cpu.scala 46:20]
  reg [31:0] DMemory_470; // @[cpu.scala 46:20]
  reg [31:0] DMemory_471; // @[cpu.scala 46:20]
  reg [31:0] DMemory_472; // @[cpu.scala 46:20]
  reg [31:0] DMemory_473; // @[cpu.scala 46:20]
  reg [31:0] DMemory_474; // @[cpu.scala 46:20]
  reg [31:0] DMemory_475; // @[cpu.scala 46:20]
  reg [31:0] DMemory_476; // @[cpu.scala 46:20]
  reg [31:0] DMemory_477; // @[cpu.scala 46:20]
  reg [31:0] DMemory_478; // @[cpu.scala 46:20]
  reg [31:0] DMemory_479; // @[cpu.scala 46:20]
  reg [31:0] DMemory_480; // @[cpu.scala 46:20]
  reg [31:0] DMemory_481; // @[cpu.scala 46:20]
  reg [31:0] DMemory_482; // @[cpu.scala 46:20]
  reg [31:0] DMemory_483; // @[cpu.scala 46:20]
  reg [31:0] DMemory_484; // @[cpu.scala 46:20]
  reg [31:0] DMemory_485; // @[cpu.scala 46:20]
  reg [31:0] DMemory_486; // @[cpu.scala 46:20]
  reg [31:0] DMemory_487; // @[cpu.scala 46:20]
  reg [31:0] DMemory_488; // @[cpu.scala 46:20]
  reg [31:0] DMemory_489; // @[cpu.scala 46:20]
  reg [31:0] DMemory_490; // @[cpu.scala 46:20]
  reg [31:0] DMemory_491; // @[cpu.scala 46:20]
  reg [31:0] DMemory_492; // @[cpu.scala 46:20]
  reg [31:0] DMemory_493; // @[cpu.scala 46:20]
  reg [31:0] DMemory_494; // @[cpu.scala 46:20]
  reg [31:0] DMemory_495; // @[cpu.scala 46:20]
  reg [31:0] DMemory_496; // @[cpu.scala 46:20]
  reg [31:0] DMemory_497; // @[cpu.scala 46:20]
  reg [31:0] DMemory_498; // @[cpu.scala 46:20]
  reg [31:0] DMemory_499; // @[cpu.scala 46:20]
  reg [31:0] DMemory_500; // @[cpu.scala 46:20]
  reg [31:0] DMemory_501; // @[cpu.scala 46:20]
  reg [31:0] DMemory_502; // @[cpu.scala 46:20]
  reg [31:0] DMemory_503; // @[cpu.scala 46:20]
  reg [31:0] DMemory_504; // @[cpu.scala 46:20]
  reg [31:0] DMemory_505; // @[cpu.scala 46:20]
  reg [31:0] DMemory_506; // @[cpu.scala 46:20]
  reg [31:0] DMemory_507; // @[cpu.scala 46:20]
  reg [31:0] DMemory_508; // @[cpu.scala 46:20]
  reg [31:0] DMemory_509; // @[cpu.scala 46:20]
  reg [31:0] DMemory_510; // @[cpu.scala 46:20]
  reg [31:0] DMemory_511; // @[cpu.scala 46:20]
  reg [31:0] DMemory_512; // @[cpu.scala 46:20]
  reg [31:0] DMemory_513; // @[cpu.scala 46:20]
  reg [31:0] DMemory_514; // @[cpu.scala 46:20]
  reg [31:0] DMemory_515; // @[cpu.scala 46:20]
  reg [31:0] DMemory_516; // @[cpu.scala 46:20]
  reg [31:0] DMemory_517; // @[cpu.scala 46:20]
  reg [31:0] DMemory_518; // @[cpu.scala 46:20]
  reg [31:0] DMemory_519; // @[cpu.scala 46:20]
  reg [31:0] DMemory_520; // @[cpu.scala 46:20]
  reg [31:0] DMemory_521; // @[cpu.scala 46:20]
  reg [31:0] DMemory_522; // @[cpu.scala 46:20]
  reg [31:0] DMemory_523; // @[cpu.scala 46:20]
  reg [31:0] DMemory_524; // @[cpu.scala 46:20]
  reg [31:0] DMemory_525; // @[cpu.scala 46:20]
  reg [31:0] DMemory_526; // @[cpu.scala 46:20]
  reg [31:0] DMemory_527; // @[cpu.scala 46:20]
  reg [31:0] DMemory_528; // @[cpu.scala 46:20]
  reg [31:0] DMemory_529; // @[cpu.scala 46:20]
  reg [31:0] DMemory_530; // @[cpu.scala 46:20]
  reg [31:0] DMemory_531; // @[cpu.scala 46:20]
  reg [31:0] DMemory_532; // @[cpu.scala 46:20]
  reg [31:0] DMemory_533; // @[cpu.scala 46:20]
  reg [31:0] DMemory_534; // @[cpu.scala 46:20]
  reg [31:0] DMemory_535; // @[cpu.scala 46:20]
  reg [31:0] DMemory_536; // @[cpu.scala 46:20]
  reg [31:0] DMemory_537; // @[cpu.scala 46:20]
  reg [31:0] DMemory_538; // @[cpu.scala 46:20]
  reg [31:0] DMemory_539; // @[cpu.scala 46:20]
  reg [31:0] DMemory_540; // @[cpu.scala 46:20]
  reg [31:0] DMemory_541; // @[cpu.scala 46:20]
  reg [31:0] DMemory_542; // @[cpu.scala 46:20]
  reg [31:0] DMemory_543; // @[cpu.scala 46:20]
  reg [31:0] DMemory_544; // @[cpu.scala 46:20]
  reg [31:0] DMemory_545; // @[cpu.scala 46:20]
  reg [31:0] DMemory_546; // @[cpu.scala 46:20]
  reg [31:0] DMemory_547; // @[cpu.scala 46:20]
  reg [31:0] DMemory_548; // @[cpu.scala 46:20]
  reg [31:0] DMemory_549; // @[cpu.scala 46:20]
  reg [31:0] DMemory_550; // @[cpu.scala 46:20]
  reg [31:0] DMemory_551; // @[cpu.scala 46:20]
  reg [31:0] DMemory_552; // @[cpu.scala 46:20]
  reg [31:0] DMemory_553; // @[cpu.scala 46:20]
  reg [31:0] DMemory_554; // @[cpu.scala 46:20]
  reg [31:0] DMemory_555; // @[cpu.scala 46:20]
  reg [31:0] DMemory_556; // @[cpu.scala 46:20]
  reg [31:0] DMemory_557; // @[cpu.scala 46:20]
  reg [31:0] DMemory_558; // @[cpu.scala 46:20]
  reg [31:0] DMemory_559; // @[cpu.scala 46:20]
  reg [31:0] DMemory_560; // @[cpu.scala 46:20]
  reg [31:0] DMemory_561; // @[cpu.scala 46:20]
  reg [31:0] DMemory_562; // @[cpu.scala 46:20]
  reg [31:0] DMemory_563; // @[cpu.scala 46:20]
  reg [31:0] DMemory_564; // @[cpu.scala 46:20]
  reg [31:0] DMemory_565; // @[cpu.scala 46:20]
  reg [31:0] DMemory_566; // @[cpu.scala 46:20]
  reg [31:0] DMemory_567; // @[cpu.scala 46:20]
  reg [31:0] DMemory_568; // @[cpu.scala 46:20]
  reg [31:0] DMemory_569; // @[cpu.scala 46:20]
  reg [31:0] DMemory_570; // @[cpu.scala 46:20]
  reg [31:0] DMemory_571; // @[cpu.scala 46:20]
  reg [31:0] DMemory_572; // @[cpu.scala 46:20]
  reg [31:0] DMemory_573; // @[cpu.scala 46:20]
  reg [31:0] DMemory_574; // @[cpu.scala 46:20]
  reg [31:0] DMemory_575; // @[cpu.scala 46:20]
  reg [31:0] DMemory_576; // @[cpu.scala 46:20]
  reg [31:0] DMemory_577; // @[cpu.scala 46:20]
  reg [31:0] DMemory_578; // @[cpu.scala 46:20]
  reg [31:0] DMemory_579; // @[cpu.scala 46:20]
  reg [31:0] DMemory_580; // @[cpu.scala 46:20]
  reg [31:0] DMemory_581; // @[cpu.scala 46:20]
  reg [31:0] DMemory_582; // @[cpu.scala 46:20]
  reg [31:0] DMemory_583; // @[cpu.scala 46:20]
  reg [31:0] DMemory_584; // @[cpu.scala 46:20]
  reg [31:0] DMemory_585; // @[cpu.scala 46:20]
  reg [31:0] DMemory_586; // @[cpu.scala 46:20]
  reg [31:0] DMemory_587; // @[cpu.scala 46:20]
  reg [31:0] DMemory_588; // @[cpu.scala 46:20]
  reg [31:0] DMemory_589; // @[cpu.scala 46:20]
  reg [31:0] DMemory_590; // @[cpu.scala 46:20]
  reg [31:0] DMemory_591; // @[cpu.scala 46:20]
  reg [31:0] DMemory_592; // @[cpu.scala 46:20]
  reg [31:0] DMemory_593; // @[cpu.scala 46:20]
  reg [31:0] DMemory_594; // @[cpu.scala 46:20]
  reg [31:0] DMemory_595; // @[cpu.scala 46:20]
  reg [31:0] DMemory_596; // @[cpu.scala 46:20]
  reg [31:0] DMemory_597; // @[cpu.scala 46:20]
  reg [31:0] DMemory_598; // @[cpu.scala 46:20]
  reg [31:0] DMemory_599; // @[cpu.scala 46:20]
  reg [31:0] DMemory_600; // @[cpu.scala 46:20]
  reg [31:0] DMemory_601; // @[cpu.scala 46:20]
  reg [31:0] DMemory_602; // @[cpu.scala 46:20]
  reg [31:0] DMemory_603; // @[cpu.scala 46:20]
  reg [31:0] DMemory_604; // @[cpu.scala 46:20]
  reg [31:0] DMemory_605; // @[cpu.scala 46:20]
  reg [31:0] DMemory_606; // @[cpu.scala 46:20]
  reg [31:0] DMemory_607; // @[cpu.scala 46:20]
  reg [31:0] DMemory_608; // @[cpu.scala 46:20]
  reg [31:0] DMemory_609; // @[cpu.scala 46:20]
  reg [31:0] DMemory_610; // @[cpu.scala 46:20]
  reg [31:0] DMemory_611; // @[cpu.scala 46:20]
  reg [31:0] DMemory_612; // @[cpu.scala 46:20]
  reg [31:0] DMemory_613; // @[cpu.scala 46:20]
  reg [31:0] DMemory_614; // @[cpu.scala 46:20]
  reg [31:0] DMemory_615; // @[cpu.scala 46:20]
  reg [31:0] DMemory_616; // @[cpu.scala 46:20]
  reg [31:0] DMemory_617; // @[cpu.scala 46:20]
  reg [31:0] DMemory_618; // @[cpu.scala 46:20]
  reg [31:0] DMemory_619; // @[cpu.scala 46:20]
  reg [31:0] DMemory_620; // @[cpu.scala 46:20]
  reg [31:0] DMemory_621; // @[cpu.scala 46:20]
  reg [31:0] DMemory_622; // @[cpu.scala 46:20]
  reg [31:0] DMemory_623; // @[cpu.scala 46:20]
  reg [31:0] DMemory_624; // @[cpu.scala 46:20]
  reg [31:0] DMemory_625; // @[cpu.scala 46:20]
  reg [31:0] DMemory_626; // @[cpu.scala 46:20]
  reg [31:0] DMemory_627; // @[cpu.scala 46:20]
  reg [31:0] DMemory_628; // @[cpu.scala 46:20]
  reg [31:0] DMemory_629; // @[cpu.scala 46:20]
  reg [31:0] DMemory_630; // @[cpu.scala 46:20]
  reg [31:0] DMemory_631; // @[cpu.scala 46:20]
  reg [31:0] DMemory_632; // @[cpu.scala 46:20]
  reg [31:0] DMemory_633; // @[cpu.scala 46:20]
  reg [31:0] DMemory_634; // @[cpu.scala 46:20]
  reg [31:0] DMemory_635; // @[cpu.scala 46:20]
  reg [31:0] DMemory_636; // @[cpu.scala 46:20]
  reg [31:0] DMemory_637; // @[cpu.scala 46:20]
  reg [31:0] DMemory_638; // @[cpu.scala 46:20]
  reg [31:0] DMemory_639; // @[cpu.scala 46:20]
  reg [31:0] DMemory_640; // @[cpu.scala 46:20]
  reg [31:0] DMemory_641; // @[cpu.scala 46:20]
  reg [31:0] DMemory_642; // @[cpu.scala 46:20]
  reg [31:0] DMemory_643; // @[cpu.scala 46:20]
  reg [31:0] DMemory_644; // @[cpu.scala 46:20]
  reg [31:0] DMemory_645; // @[cpu.scala 46:20]
  reg [31:0] DMemory_646; // @[cpu.scala 46:20]
  reg [31:0] DMemory_647; // @[cpu.scala 46:20]
  reg [31:0] DMemory_648; // @[cpu.scala 46:20]
  reg [31:0] DMemory_649; // @[cpu.scala 46:20]
  reg [31:0] DMemory_650; // @[cpu.scala 46:20]
  reg [31:0] DMemory_651; // @[cpu.scala 46:20]
  reg [31:0] DMemory_652; // @[cpu.scala 46:20]
  reg [31:0] DMemory_653; // @[cpu.scala 46:20]
  reg [31:0] DMemory_654; // @[cpu.scala 46:20]
  reg [31:0] DMemory_655; // @[cpu.scala 46:20]
  reg [31:0] DMemory_656; // @[cpu.scala 46:20]
  reg [31:0] DMemory_657; // @[cpu.scala 46:20]
  reg [31:0] DMemory_658; // @[cpu.scala 46:20]
  reg [31:0] DMemory_659; // @[cpu.scala 46:20]
  reg [31:0] DMemory_660; // @[cpu.scala 46:20]
  reg [31:0] DMemory_661; // @[cpu.scala 46:20]
  reg [31:0] DMemory_662; // @[cpu.scala 46:20]
  reg [31:0] DMemory_663; // @[cpu.scala 46:20]
  reg [31:0] DMemory_664; // @[cpu.scala 46:20]
  reg [31:0] DMemory_665; // @[cpu.scala 46:20]
  reg [31:0] DMemory_666; // @[cpu.scala 46:20]
  reg [31:0] DMemory_667; // @[cpu.scala 46:20]
  reg [31:0] DMemory_668; // @[cpu.scala 46:20]
  reg [31:0] DMemory_669; // @[cpu.scala 46:20]
  reg [31:0] DMemory_670; // @[cpu.scala 46:20]
  reg [31:0] DMemory_671; // @[cpu.scala 46:20]
  reg [31:0] DMemory_672; // @[cpu.scala 46:20]
  reg [31:0] DMemory_673; // @[cpu.scala 46:20]
  reg [31:0] DMemory_674; // @[cpu.scala 46:20]
  reg [31:0] DMemory_675; // @[cpu.scala 46:20]
  reg [31:0] DMemory_676; // @[cpu.scala 46:20]
  reg [31:0] DMemory_677; // @[cpu.scala 46:20]
  reg [31:0] DMemory_678; // @[cpu.scala 46:20]
  reg [31:0] DMemory_679; // @[cpu.scala 46:20]
  reg [31:0] DMemory_680; // @[cpu.scala 46:20]
  reg [31:0] DMemory_681; // @[cpu.scala 46:20]
  reg [31:0] DMemory_682; // @[cpu.scala 46:20]
  reg [31:0] DMemory_683; // @[cpu.scala 46:20]
  reg [31:0] DMemory_684; // @[cpu.scala 46:20]
  reg [31:0] DMemory_685; // @[cpu.scala 46:20]
  reg [31:0] DMemory_686; // @[cpu.scala 46:20]
  reg [31:0] DMemory_687; // @[cpu.scala 46:20]
  reg [31:0] DMemory_688; // @[cpu.scala 46:20]
  reg [31:0] DMemory_689; // @[cpu.scala 46:20]
  reg [31:0] DMemory_690; // @[cpu.scala 46:20]
  reg [31:0] DMemory_691; // @[cpu.scala 46:20]
  reg [31:0] DMemory_692; // @[cpu.scala 46:20]
  reg [31:0] DMemory_693; // @[cpu.scala 46:20]
  reg [31:0] DMemory_694; // @[cpu.scala 46:20]
  reg [31:0] DMemory_695; // @[cpu.scala 46:20]
  reg [31:0] DMemory_696; // @[cpu.scala 46:20]
  reg [31:0] DMemory_697; // @[cpu.scala 46:20]
  reg [31:0] DMemory_698; // @[cpu.scala 46:20]
  reg [31:0] DMemory_699; // @[cpu.scala 46:20]
  reg [31:0] DMemory_700; // @[cpu.scala 46:20]
  reg [31:0] DMemory_701; // @[cpu.scala 46:20]
  reg [31:0] DMemory_702; // @[cpu.scala 46:20]
  reg [31:0] DMemory_703; // @[cpu.scala 46:20]
  reg [31:0] DMemory_704; // @[cpu.scala 46:20]
  reg [31:0] DMemory_705; // @[cpu.scala 46:20]
  reg [31:0] DMemory_706; // @[cpu.scala 46:20]
  reg [31:0] DMemory_707; // @[cpu.scala 46:20]
  reg [31:0] DMemory_708; // @[cpu.scala 46:20]
  reg [31:0] DMemory_709; // @[cpu.scala 46:20]
  reg [31:0] DMemory_710; // @[cpu.scala 46:20]
  reg [31:0] DMemory_711; // @[cpu.scala 46:20]
  reg [31:0] DMemory_712; // @[cpu.scala 46:20]
  reg [31:0] DMemory_713; // @[cpu.scala 46:20]
  reg [31:0] DMemory_714; // @[cpu.scala 46:20]
  reg [31:0] DMemory_715; // @[cpu.scala 46:20]
  reg [31:0] DMemory_716; // @[cpu.scala 46:20]
  reg [31:0] DMemory_717; // @[cpu.scala 46:20]
  reg [31:0] DMemory_718; // @[cpu.scala 46:20]
  reg [31:0] DMemory_719; // @[cpu.scala 46:20]
  reg [31:0] DMemory_720; // @[cpu.scala 46:20]
  reg [31:0] DMemory_721; // @[cpu.scala 46:20]
  reg [31:0] DMemory_722; // @[cpu.scala 46:20]
  reg [31:0] DMemory_723; // @[cpu.scala 46:20]
  reg [31:0] DMemory_724; // @[cpu.scala 46:20]
  reg [31:0] DMemory_725; // @[cpu.scala 46:20]
  reg [31:0] DMemory_726; // @[cpu.scala 46:20]
  reg [31:0] DMemory_727; // @[cpu.scala 46:20]
  reg [31:0] DMemory_728; // @[cpu.scala 46:20]
  reg [31:0] DMemory_729; // @[cpu.scala 46:20]
  reg [31:0] DMemory_730; // @[cpu.scala 46:20]
  reg [31:0] DMemory_731; // @[cpu.scala 46:20]
  reg [31:0] DMemory_732; // @[cpu.scala 46:20]
  reg [31:0] DMemory_733; // @[cpu.scala 46:20]
  reg [31:0] DMemory_734; // @[cpu.scala 46:20]
  reg [31:0] DMemory_735; // @[cpu.scala 46:20]
  reg [31:0] DMemory_736; // @[cpu.scala 46:20]
  reg [31:0] DMemory_737; // @[cpu.scala 46:20]
  reg [31:0] DMemory_738; // @[cpu.scala 46:20]
  reg [31:0] DMemory_739; // @[cpu.scala 46:20]
  reg [31:0] DMemory_740; // @[cpu.scala 46:20]
  reg [31:0] DMemory_741; // @[cpu.scala 46:20]
  reg [31:0] DMemory_742; // @[cpu.scala 46:20]
  reg [31:0] DMemory_743; // @[cpu.scala 46:20]
  reg [31:0] DMemory_744; // @[cpu.scala 46:20]
  reg [31:0] DMemory_745; // @[cpu.scala 46:20]
  reg [31:0] DMemory_746; // @[cpu.scala 46:20]
  reg [31:0] DMemory_747; // @[cpu.scala 46:20]
  reg [31:0] DMemory_748; // @[cpu.scala 46:20]
  reg [31:0] DMemory_749; // @[cpu.scala 46:20]
  reg [31:0] DMemory_750; // @[cpu.scala 46:20]
  reg [31:0] DMemory_751; // @[cpu.scala 46:20]
  reg [31:0] DMemory_752; // @[cpu.scala 46:20]
  reg [31:0] DMemory_753; // @[cpu.scala 46:20]
  reg [31:0] DMemory_754; // @[cpu.scala 46:20]
  reg [31:0] DMemory_755; // @[cpu.scala 46:20]
  reg [31:0] DMemory_756; // @[cpu.scala 46:20]
  reg [31:0] DMemory_757; // @[cpu.scala 46:20]
  reg [31:0] DMemory_758; // @[cpu.scala 46:20]
  reg [31:0] DMemory_759; // @[cpu.scala 46:20]
  reg [31:0] DMemory_760; // @[cpu.scala 46:20]
  reg [31:0] DMemory_761; // @[cpu.scala 46:20]
  reg [31:0] DMemory_762; // @[cpu.scala 46:20]
  reg [31:0] DMemory_763; // @[cpu.scala 46:20]
  reg [31:0] DMemory_764; // @[cpu.scala 46:20]
  reg [31:0] DMemory_765; // @[cpu.scala 46:20]
  reg [31:0] DMemory_766; // @[cpu.scala 46:20]
  reg [31:0] DMemory_767; // @[cpu.scala 46:20]
  reg [31:0] DMemory_768; // @[cpu.scala 46:20]
  reg [31:0] DMemory_769; // @[cpu.scala 46:20]
  reg [31:0] DMemory_770; // @[cpu.scala 46:20]
  reg [31:0] DMemory_771; // @[cpu.scala 46:20]
  reg [31:0] DMemory_772; // @[cpu.scala 46:20]
  reg [31:0] DMemory_773; // @[cpu.scala 46:20]
  reg [31:0] DMemory_774; // @[cpu.scala 46:20]
  reg [31:0] DMemory_775; // @[cpu.scala 46:20]
  reg [31:0] DMemory_776; // @[cpu.scala 46:20]
  reg [31:0] DMemory_777; // @[cpu.scala 46:20]
  reg [31:0] DMemory_778; // @[cpu.scala 46:20]
  reg [31:0] DMemory_779; // @[cpu.scala 46:20]
  reg [31:0] DMemory_780; // @[cpu.scala 46:20]
  reg [31:0] DMemory_781; // @[cpu.scala 46:20]
  reg [31:0] DMemory_782; // @[cpu.scala 46:20]
  reg [31:0] DMemory_783; // @[cpu.scala 46:20]
  reg [31:0] DMemory_784; // @[cpu.scala 46:20]
  reg [31:0] DMemory_785; // @[cpu.scala 46:20]
  reg [31:0] DMemory_786; // @[cpu.scala 46:20]
  reg [31:0] DMemory_787; // @[cpu.scala 46:20]
  reg [31:0] DMemory_788; // @[cpu.scala 46:20]
  reg [31:0] DMemory_789; // @[cpu.scala 46:20]
  reg [31:0] DMemory_790; // @[cpu.scala 46:20]
  reg [31:0] DMemory_791; // @[cpu.scala 46:20]
  reg [31:0] DMemory_792; // @[cpu.scala 46:20]
  reg [31:0] DMemory_793; // @[cpu.scala 46:20]
  reg [31:0] DMemory_794; // @[cpu.scala 46:20]
  reg [31:0] DMemory_795; // @[cpu.scala 46:20]
  reg [31:0] DMemory_796; // @[cpu.scala 46:20]
  reg [31:0] DMemory_797; // @[cpu.scala 46:20]
  reg [31:0] DMemory_798; // @[cpu.scala 46:20]
  reg [31:0] DMemory_799; // @[cpu.scala 46:20]
  reg [31:0] DMemory_800; // @[cpu.scala 46:20]
  reg [31:0] DMemory_801; // @[cpu.scala 46:20]
  reg [31:0] DMemory_802; // @[cpu.scala 46:20]
  reg [31:0] DMemory_803; // @[cpu.scala 46:20]
  reg [31:0] DMemory_804; // @[cpu.scala 46:20]
  reg [31:0] DMemory_805; // @[cpu.scala 46:20]
  reg [31:0] DMemory_806; // @[cpu.scala 46:20]
  reg [31:0] DMemory_807; // @[cpu.scala 46:20]
  reg [31:0] DMemory_808; // @[cpu.scala 46:20]
  reg [31:0] DMemory_809; // @[cpu.scala 46:20]
  reg [31:0] DMemory_810; // @[cpu.scala 46:20]
  reg [31:0] DMemory_811; // @[cpu.scala 46:20]
  reg [31:0] DMemory_812; // @[cpu.scala 46:20]
  reg [31:0] DMemory_813; // @[cpu.scala 46:20]
  reg [31:0] DMemory_814; // @[cpu.scala 46:20]
  reg [31:0] DMemory_815; // @[cpu.scala 46:20]
  reg [31:0] DMemory_816; // @[cpu.scala 46:20]
  reg [31:0] DMemory_817; // @[cpu.scala 46:20]
  reg [31:0] DMemory_818; // @[cpu.scala 46:20]
  reg [31:0] DMemory_819; // @[cpu.scala 46:20]
  reg [31:0] DMemory_820; // @[cpu.scala 46:20]
  reg [31:0] DMemory_821; // @[cpu.scala 46:20]
  reg [31:0] DMemory_822; // @[cpu.scala 46:20]
  reg [31:0] DMemory_823; // @[cpu.scala 46:20]
  reg [31:0] DMemory_824; // @[cpu.scala 46:20]
  reg [31:0] DMemory_825; // @[cpu.scala 46:20]
  reg [31:0] DMemory_826; // @[cpu.scala 46:20]
  reg [31:0] DMemory_827; // @[cpu.scala 46:20]
  reg [31:0] DMemory_828; // @[cpu.scala 46:20]
  reg [31:0] DMemory_829; // @[cpu.scala 46:20]
  reg [31:0] DMemory_830; // @[cpu.scala 46:20]
  reg [31:0] DMemory_831; // @[cpu.scala 46:20]
  reg [31:0] DMemory_832; // @[cpu.scala 46:20]
  reg [31:0] DMemory_833; // @[cpu.scala 46:20]
  reg [31:0] DMemory_834; // @[cpu.scala 46:20]
  reg [31:0] DMemory_835; // @[cpu.scala 46:20]
  reg [31:0] DMemory_836; // @[cpu.scala 46:20]
  reg [31:0] DMemory_837; // @[cpu.scala 46:20]
  reg [31:0] DMemory_838; // @[cpu.scala 46:20]
  reg [31:0] DMemory_839; // @[cpu.scala 46:20]
  reg [31:0] DMemory_840; // @[cpu.scala 46:20]
  reg [31:0] DMemory_841; // @[cpu.scala 46:20]
  reg [31:0] DMemory_842; // @[cpu.scala 46:20]
  reg [31:0] DMemory_843; // @[cpu.scala 46:20]
  reg [31:0] DMemory_844; // @[cpu.scala 46:20]
  reg [31:0] DMemory_845; // @[cpu.scala 46:20]
  reg [31:0] DMemory_846; // @[cpu.scala 46:20]
  reg [31:0] DMemory_847; // @[cpu.scala 46:20]
  reg [31:0] DMemory_848; // @[cpu.scala 46:20]
  reg [31:0] DMemory_849; // @[cpu.scala 46:20]
  reg [31:0] DMemory_850; // @[cpu.scala 46:20]
  reg [31:0] DMemory_851; // @[cpu.scala 46:20]
  reg [31:0] DMemory_852; // @[cpu.scala 46:20]
  reg [31:0] DMemory_853; // @[cpu.scala 46:20]
  reg [31:0] DMemory_854; // @[cpu.scala 46:20]
  reg [31:0] DMemory_855; // @[cpu.scala 46:20]
  reg [31:0] DMemory_856; // @[cpu.scala 46:20]
  reg [31:0] DMemory_857; // @[cpu.scala 46:20]
  reg [31:0] DMemory_858; // @[cpu.scala 46:20]
  reg [31:0] DMemory_859; // @[cpu.scala 46:20]
  reg [31:0] DMemory_860; // @[cpu.scala 46:20]
  reg [31:0] DMemory_861; // @[cpu.scala 46:20]
  reg [31:0] DMemory_862; // @[cpu.scala 46:20]
  reg [31:0] DMemory_863; // @[cpu.scala 46:20]
  reg [31:0] DMemory_864; // @[cpu.scala 46:20]
  reg [31:0] DMemory_865; // @[cpu.scala 46:20]
  reg [31:0] DMemory_866; // @[cpu.scala 46:20]
  reg [31:0] DMemory_867; // @[cpu.scala 46:20]
  reg [31:0] DMemory_868; // @[cpu.scala 46:20]
  reg [31:0] DMemory_869; // @[cpu.scala 46:20]
  reg [31:0] DMemory_870; // @[cpu.scala 46:20]
  reg [31:0] DMemory_871; // @[cpu.scala 46:20]
  reg [31:0] DMemory_872; // @[cpu.scala 46:20]
  reg [31:0] DMemory_873; // @[cpu.scala 46:20]
  reg [31:0] DMemory_874; // @[cpu.scala 46:20]
  reg [31:0] DMemory_875; // @[cpu.scala 46:20]
  reg [31:0] DMemory_876; // @[cpu.scala 46:20]
  reg [31:0] DMemory_877; // @[cpu.scala 46:20]
  reg [31:0] DMemory_878; // @[cpu.scala 46:20]
  reg [31:0] DMemory_879; // @[cpu.scala 46:20]
  reg [31:0] DMemory_880; // @[cpu.scala 46:20]
  reg [31:0] DMemory_881; // @[cpu.scala 46:20]
  reg [31:0] DMemory_882; // @[cpu.scala 46:20]
  reg [31:0] DMemory_883; // @[cpu.scala 46:20]
  reg [31:0] DMemory_884; // @[cpu.scala 46:20]
  reg [31:0] DMemory_885; // @[cpu.scala 46:20]
  reg [31:0] DMemory_886; // @[cpu.scala 46:20]
  reg [31:0] DMemory_887; // @[cpu.scala 46:20]
  reg [31:0] DMemory_888; // @[cpu.scala 46:20]
  reg [31:0] DMemory_889; // @[cpu.scala 46:20]
  reg [31:0] DMemory_890; // @[cpu.scala 46:20]
  reg [31:0] DMemory_891; // @[cpu.scala 46:20]
  reg [31:0] DMemory_892; // @[cpu.scala 46:20]
  reg [31:0] DMemory_893; // @[cpu.scala 46:20]
  reg [31:0] DMemory_894; // @[cpu.scala 46:20]
  reg [31:0] DMemory_895; // @[cpu.scala 46:20]
  reg [31:0] DMemory_896; // @[cpu.scala 46:20]
  reg [31:0] DMemory_897; // @[cpu.scala 46:20]
  reg [31:0] DMemory_898; // @[cpu.scala 46:20]
  reg [31:0] DMemory_899; // @[cpu.scala 46:20]
  reg [31:0] DMemory_900; // @[cpu.scala 46:20]
  reg [31:0] DMemory_901; // @[cpu.scala 46:20]
  reg [31:0] DMemory_902; // @[cpu.scala 46:20]
  reg [31:0] DMemory_903; // @[cpu.scala 46:20]
  reg [31:0] DMemory_904; // @[cpu.scala 46:20]
  reg [31:0] DMemory_905; // @[cpu.scala 46:20]
  reg [31:0] DMemory_906; // @[cpu.scala 46:20]
  reg [31:0] DMemory_907; // @[cpu.scala 46:20]
  reg [31:0] DMemory_908; // @[cpu.scala 46:20]
  reg [31:0] DMemory_909; // @[cpu.scala 46:20]
  reg [31:0] DMemory_910; // @[cpu.scala 46:20]
  reg [31:0] DMemory_911; // @[cpu.scala 46:20]
  reg [31:0] DMemory_912; // @[cpu.scala 46:20]
  reg [31:0] DMemory_913; // @[cpu.scala 46:20]
  reg [31:0] DMemory_914; // @[cpu.scala 46:20]
  reg [31:0] DMemory_915; // @[cpu.scala 46:20]
  reg [31:0] DMemory_916; // @[cpu.scala 46:20]
  reg [31:0] DMemory_917; // @[cpu.scala 46:20]
  reg [31:0] DMemory_918; // @[cpu.scala 46:20]
  reg [31:0] DMemory_919; // @[cpu.scala 46:20]
  reg [31:0] DMemory_920; // @[cpu.scala 46:20]
  reg [31:0] DMemory_921; // @[cpu.scala 46:20]
  reg [31:0] DMemory_922; // @[cpu.scala 46:20]
  reg [31:0] DMemory_923; // @[cpu.scala 46:20]
  reg [31:0] DMemory_924; // @[cpu.scala 46:20]
  reg [31:0] DMemory_925; // @[cpu.scala 46:20]
  reg [31:0] DMemory_926; // @[cpu.scala 46:20]
  reg [31:0] DMemory_927; // @[cpu.scala 46:20]
  reg [31:0] DMemory_928; // @[cpu.scala 46:20]
  reg [31:0] DMemory_929; // @[cpu.scala 46:20]
  reg [31:0] DMemory_930; // @[cpu.scala 46:20]
  reg [31:0] DMemory_931; // @[cpu.scala 46:20]
  reg [31:0] DMemory_932; // @[cpu.scala 46:20]
  reg [31:0] DMemory_933; // @[cpu.scala 46:20]
  reg [31:0] DMemory_934; // @[cpu.scala 46:20]
  reg [31:0] DMemory_935; // @[cpu.scala 46:20]
  reg [31:0] DMemory_936; // @[cpu.scala 46:20]
  reg [31:0] DMemory_937; // @[cpu.scala 46:20]
  reg [31:0] DMemory_938; // @[cpu.scala 46:20]
  reg [31:0] DMemory_939; // @[cpu.scala 46:20]
  reg [31:0] DMemory_940; // @[cpu.scala 46:20]
  reg [31:0] DMemory_941; // @[cpu.scala 46:20]
  reg [31:0] DMemory_942; // @[cpu.scala 46:20]
  reg [31:0] DMemory_943; // @[cpu.scala 46:20]
  reg [31:0] DMemory_944; // @[cpu.scala 46:20]
  reg [31:0] DMemory_945; // @[cpu.scala 46:20]
  reg [31:0] DMemory_946; // @[cpu.scala 46:20]
  reg [31:0] DMemory_947; // @[cpu.scala 46:20]
  reg [31:0] DMemory_948; // @[cpu.scala 46:20]
  reg [31:0] DMemory_949; // @[cpu.scala 46:20]
  reg [31:0] DMemory_950; // @[cpu.scala 46:20]
  reg [31:0] DMemory_951; // @[cpu.scala 46:20]
  reg [31:0] DMemory_952; // @[cpu.scala 46:20]
  reg [31:0] DMemory_953; // @[cpu.scala 46:20]
  reg [31:0] DMemory_954; // @[cpu.scala 46:20]
  reg [31:0] DMemory_955; // @[cpu.scala 46:20]
  reg [31:0] DMemory_956; // @[cpu.scala 46:20]
  reg [31:0] DMemory_957; // @[cpu.scala 46:20]
  reg [31:0] DMemory_958; // @[cpu.scala 46:20]
  reg [31:0] DMemory_959; // @[cpu.scala 46:20]
  reg [31:0] DMemory_960; // @[cpu.scala 46:20]
  reg [31:0] DMemory_961; // @[cpu.scala 46:20]
  reg [31:0] DMemory_962; // @[cpu.scala 46:20]
  reg [31:0] DMemory_963; // @[cpu.scala 46:20]
  reg [31:0] DMemory_964; // @[cpu.scala 46:20]
  reg [31:0] DMemory_965; // @[cpu.scala 46:20]
  reg [31:0] DMemory_966; // @[cpu.scala 46:20]
  reg [31:0] DMemory_967; // @[cpu.scala 46:20]
  reg [31:0] DMemory_968; // @[cpu.scala 46:20]
  reg [31:0] DMemory_969; // @[cpu.scala 46:20]
  reg [31:0] DMemory_970; // @[cpu.scala 46:20]
  reg [31:0] DMemory_971; // @[cpu.scala 46:20]
  reg [31:0] DMemory_972; // @[cpu.scala 46:20]
  reg [31:0] DMemory_973; // @[cpu.scala 46:20]
  reg [31:0] DMemory_974; // @[cpu.scala 46:20]
  reg [31:0] DMemory_975; // @[cpu.scala 46:20]
  reg [31:0] DMemory_976; // @[cpu.scala 46:20]
  reg [31:0] DMemory_977; // @[cpu.scala 46:20]
  reg [31:0] DMemory_978; // @[cpu.scala 46:20]
  reg [31:0] DMemory_979; // @[cpu.scala 46:20]
  reg [31:0] DMemory_980; // @[cpu.scala 46:20]
  reg [31:0] DMemory_981; // @[cpu.scala 46:20]
  reg [31:0] DMemory_982; // @[cpu.scala 46:20]
  reg [31:0] DMemory_983; // @[cpu.scala 46:20]
  reg [31:0] DMemory_984; // @[cpu.scala 46:20]
  reg [31:0] DMemory_985; // @[cpu.scala 46:20]
  reg [31:0] DMemory_986; // @[cpu.scala 46:20]
  reg [31:0] DMemory_987; // @[cpu.scala 46:20]
  reg [31:0] DMemory_988; // @[cpu.scala 46:20]
  reg [31:0] DMemory_989; // @[cpu.scala 46:20]
  reg [31:0] DMemory_990; // @[cpu.scala 46:20]
  reg [31:0] DMemory_991; // @[cpu.scala 46:20]
  reg [31:0] DMemory_992; // @[cpu.scala 46:20]
  reg [31:0] DMemory_993; // @[cpu.scala 46:20]
  reg [31:0] DMemory_994; // @[cpu.scala 46:20]
  reg [31:0] DMemory_995; // @[cpu.scala 46:20]
  reg [31:0] DMemory_996; // @[cpu.scala 46:20]
  reg [31:0] DMemory_997; // @[cpu.scala 46:20]
  reg [31:0] DMemory_998; // @[cpu.scala 46:20]
  reg [31:0] DMemory_999; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1000; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1001; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1002; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1003; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1004; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1005; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1006; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1007; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1008; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1009; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1010; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1011; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1012; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1013; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1014; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1015; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1016; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1017; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1018; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1019; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1020; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1021; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1022; // @[cpu.scala 46:20]
  reg [31:0] DMemory_1023; // @[cpu.scala 46:20]
  reg [31:0] IMemory_0; // @[cpu.scala 47:20]
  reg [31:0] IMemory_1; // @[cpu.scala 47:20]
  reg [31:0] IMemory_2; // @[cpu.scala 47:20]
  reg [31:0] IMemory_3; // @[cpu.scala 47:20]
  reg [31:0] IMemory_4; // @[cpu.scala 47:20]
  reg [31:0] IMemory_5; // @[cpu.scala 47:20]
  reg [31:0] IMemory_6; // @[cpu.scala 47:20]
  reg [31:0] IMemory_7; // @[cpu.scala 47:20]
  reg [31:0] IFIDIR; // @[cpu.scala 48:49]
  reg [31:0] IDEXIR; // @[cpu.scala 48:49]
  reg [31:0] EXMEMIR; // @[cpu.scala 48:49]
  reg [31:0] MEMWBIR; // @[cpu.scala 48:49]
  reg [63:0] CurPC; // @[cpu.scala 51:22]
  wire [4:0] EXMEMrd = EXMEMIR[11:7]; // @[cpu.scala 85:32]
  wire [4:0] IDEXrd = IDEXIR[11:7]; // @[cpu.scala 86:30]
  wire [2:0] IFID_funct3 = IFIDIR[14:12]; // @[cpu.scala 87:29]
  wire [4:0] IFIDrs1 = io_rvfi_rst ? IFIDIR[19:15] : IFIDIR[19:15]; // @[cpu.scala 55:21 57:13 77:13]
  wire [4:0] MEMWBrd = io_rvfi_rst ? MEMWBIR[11:7] : MEMWBIR[11:7]; // @[cpu.scala 55:21 63:13 83:13]
  wire  _bypassAFromWB_T_1 = IFIDrs1 != 5'h0; // @[cpu.scala 90:41]
  wire [6:0] MEMWBop = io_rvfi_rst ? MEMWBIR[6:0] : MEMWBIR[6:0]; // @[cpu.scala 55:21 62:13 82:13]
  wire  _bypassAFromWB_T_3 = MEMWBop == 7'h33; // @[cpu.scala 90:62]
  wire  _bypassAFromWB_T_4 = MEMWBop == 7'h3; // @[cpu.scala 90:83]
  wire  _bypassAFromWB_T_5 = MEMWBop == 7'h33 | MEMWBop == 7'h3; // @[cpu.scala 90:72]
  wire  bypassAFromWB = IFIDrs1 == MEMWBrd & IFIDrs1 != 5'h0 & (MEMWBop == 7'h33 | MEMWBop == 7'h3); // @[cpu.scala 90:50]
  wire [4:0] IFIDrs2 = io_rvfi_rst ? IFIDIR[24:20] : IFIDIR[24:20]; // @[cpu.scala 55:21 58:13 78:13]
  wire  _bypassBFromWB_T_1 = IFIDrs2 != 5'h0; // @[cpu.scala 92:41]
  wire  bypassBFromWB = IFIDrs2 == MEMWBrd & IFIDrs2 != 5'h0 & _bypassAFromWB_T_5; // @[cpu.scala 92:50]
  wire  _bypassAFromMEM_T_2 = IFIDrs1 == EXMEMrd & _bypassAFromWB_T_1; // @[cpu.scala 94:29]
  wire [6:0] EXMEMop = io_rvfi_rst ? EXMEMIR[6:0] : EXMEMIR[6:0]; // @[cpu.scala 55:21 61:13 81:13]
  wire  _bypassAFromMEM_T_3 = EXMEMop == 7'h33; // @[cpu.scala 94:62]
  wire  bypassAFromMEM = IFIDrs1 == EXMEMrd & _bypassAFromWB_T_1 & EXMEMop == 7'h33; // @[cpu.scala 94:50]
  wire  _bypassBFromMEM_T_2 = IFIDrs2 == EXMEMrd & _bypassBFromWB_T_1; // @[cpu.scala 96:29]
  wire  bypassBFromMEM = IFIDrs2 == EXMEMrd & _bypassBFromWB_T_1 & _bypassAFromMEM_T_3; // @[cpu.scala 96:50]
  wire  _bypassAFromEX_T_2 = IFIDrs1 == IDEXrd & _bypassAFromWB_T_1; // @[cpu.scala 98:28]
  wire [6:0] IDEXop = io_rvfi_rst ? IDEXIR[6:0] : IDEXIR[6:0]; // @[cpu.scala 55:21 59:12 79:12]
  wire  _bypassAFromEX_T_3 = IDEXop == 7'h33; // @[cpu.scala 98:60]
  wire  bypassAFromEX = IFIDrs1 == IDEXrd & _bypassAFromWB_T_1 & IDEXop == 7'h33; // @[cpu.scala 98:49]
  wire  _bypassBFromEX_T_2 = IFIDrs2 == IDEXrd & _bypassBFromWB_T_1; // @[cpu.scala 100:28]
  wire  bypassBFromEX = IFIDrs2 == IDEXrd & _bypassBFromWB_T_1 & _bypassAFromEX_T_3; // @[cpu.scala 100:49]
  wire  _stall_T = EXMEMop == 7'h3; // @[cpu.scala 103:16]
  wire  _stall_T_8 = EXMEMop == 7'h3 & (_bypassAFromMEM_T_2 | _bypassBFromMEM_T_2); // @[cpu.scala 103:24]
  wire  _stall_T_9 = IDEXop == 7'h3; // @[cpu.scala 105:15]
  wire  _stall_T_17 = IDEXop == 7'h3 & (_bypassAFromEX_T_2 | _bypassBFromEX_T_2); // @[cpu.scala 105:23]
  wire  stall = _stall_T_8 | _stall_T_17; // @[cpu.scala 104:7]
  wire [6:0] IFIDop = io_rvfi_rst ? IFIDIR[6:0] : IFIDIR[6:0]; // @[cpu.scala 55:21 60:12 80:12]
  wire [63:0] _A_T_1 = IDEXA + IDEXB; // @[cpu.scala 146:20]
  wire [63:0] _GEN_1029 = 5'h1 == IFIDrs1 ? Regs_1 : Regs_0; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1030 = 5'h2 == IFIDrs1 ? Regs_2 : _GEN_1029; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1031 = 5'h3 == IFIDrs1 ? Regs_3 : _GEN_1030; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1032 = 5'h4 == IFIDrs1 ? Regs_4 : _GEN_1031; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1033 = 5'h5 == IFIDrs1 ? Regs_5 : _GEN_1032; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1034 = 5'h6 == IFIDrs1 ? Regs_6 : _GEN_1033; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1035 = 5'h7 == IFIDrs1 ? Regs_7 : _GEN_1034; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1036 = 5'h8 == IFIDrs1 ? Regs_8 : _GEN_1035; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1037 = 5'h9 == IFIDrs1 ? Regs_9 : _GEN_1036; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1038 = 5'ha == IFIDrs1 ? Regs_10 : _GEN_1037; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1039 = 5'hb == IFIDrs1 ? Regs_11 : _GEN_1038; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1040 = 5'hc == IFIDrs1 ? Regs_12 : _GEN_1039; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1041 = 5'hd == IFIDrs1 ? Regs_13 : _GEN_1040; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1042 = 5'he == IFIDrs1 ? Regs_14 : _GEN_1041; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1043 = 5'hf == IFIDrs1 ? Regs_15 : _GEN_1042; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1044 = 5'h10 == IFIDrs1 ? Regs_16 : _GEN_1043; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1045 = 5'h11 == IFIDrs1 ? Regs_17 : _GEN_1044; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1046 = 5'h12 == IFIDrs1 ? Regs_18 : _GEN_1045; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1047 = 5'h13 == IFIDrs1 ? Regs_19 : _GEN_1046; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1048 = 5'h14 == IFIDrs1 ? Regs_20 : _GEN_1047; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1049 = 5'h15 == IFIDrs1 ? Regs_21 : _GEN_1048; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1050 = 5'h16 == IFIDrs1 ? Regs_22 : _GEN_1049; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1051 = 5'h17 == IFIDrs1 ? Regs_23 : _GEN_1050; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1052 = 5'h18 == IFIDrs1 ? Regs_24 : _GEN_1051; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1053 = 5'h19 == IFIDrs1 ? Regs_25 : _GEN_1052; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1054 = 5'h1a == IFIDrs1 ? Regs_26 : _GEN_1053; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1055 = 5'h1b == IFIDrs1 ? Regs_27 : _GEN_1054; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1056 = 5'h1c == IFIDrs1 ? Regs_28 : _GEN_1055; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1057 = 5'h1d == IFIDrs1 ? Regs_29 : _GEN_1056; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1058 = 5'h1e == IFIDrs1 ? Regs_30 : _GEN_1057; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1059 = 5'h1f == IFIDrs1 ? Regs_31 : _GEN_1058; // @[cpu.scala 154:{15,15}]
  wire [63:0] _GEN_1061 = bypassAFromWB ? MEMWBValue : _GEN_1059; // @[cpu.scala 150:33 152:11 155:11]
  wire [63:0] _GEN_1063 = bypassAFromMEM ? EXMEMALUOut : _GEN_1061; // @[cpu.scala 147:34 149:11]
  wire [63:0] _GEN_1065 = bypassAFromEX ? _A_T_1 : _GEN_1063; // @[cpu.scala 144:27 146:11]
  wire [63:0] A = ~stall ? _GEN_1065 : 64'h0; // @[cpu.scala 117:27]
  wire [63:0] _B_T_1 = IDEXB + IDEXA; // @[cpu.scala 159:20]
  wire [63:0] _GEN_1067 = 5'h1 == IFIDrs2 ? Regs_1 : Regs_0; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1068 = 5'h2 == IFIDrs2 ? Regs_2 : _GEN_1067; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1069 = 5'h3 == IFIDrs2 ? Regs_3 : _GEN_1068; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1070 = 5'h4 == IFIDrs2 ? Regs_4 : _GEN_1069; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1071 = 5'h5 == IFIDrs2 ? Regs_5 : _GEN_1070; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1072 = 5'h6 == IFIDrs2 ? Regs_6 : _GEN_1071; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1073 = 5'h7 == IFIDrs2 ? Regs_7 : _GEN_1072; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1074 = 5'h8 == IFIDrs2 ? Regs_8 : _GEN_1073; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1075 = 5'h9 == IFIDrs2 ? Regs_9 : _GEN_1074; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1076 = 5'ha == IFIDrs2 ? Regs_10 : _GEN_1075; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1077 = 5'hb == IFIDrs2 ? Regs_11 : _GEN_1076; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1078 = 5'hc == IFIDrs2 ? Regs_12 : _GEN_1077; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1079 = 5'hd == IFIDrs2 ? Regs_13 : _GEN_1078; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1080 = 5'he == IFIDrs2 ? Regs_14 : _GEN_1079; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1081 = 5'hf == IFIDrs2 ? Regs_15 : _GEN_1080; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1082 = 5'h10 == IFIDrs2 ? Regs_16 : _GEN_1081; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1083 = 5'h11 == IFIDrs2 ? Regs_17 : _GEN_1082; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1084 = 5'h12 == IFIDrs2 ? Regs_18 : _GEN_1083; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1085 = 5'h13 == IFIDrs2 ? Regs_19 : _GEN_1084; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1086 = 5'h14 == IFIDrs2 ? Regs_20 : _GEN_1085; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1087 = 5'h15 == IFIDrs2 ? Regs_21 : _GEN_1086; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1088 = 5'h16 == IFIDrs2 ? Regs_22 : _GEN_1087; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1089 = 5'h17 == IFIDrs2 ? Regs_23 : _GEN_1088; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1090 = 5'h18 == IFIDrs2 ? Regs_24 : _GEN_1089; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1091 = 5'h19 == IFIDrs2 ? Regs_25 : _GEN_1090; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1092 = 5'h1a == IFIDrs2 ? Regs_26 : _GEN_1091; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1093 = 5'h1b == IFIDrs2 ? Regs_27 : _GEN_1092; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1094 = 5'h1c == IFIDrs2 ? Regs_28 : _GEN_1093; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1095 = 5'h1d == IFIDrs2 ? Regs_29 : _GEN_1094; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1096 = 5'h1e == IFIDrs2 ? Regs_30 : _GEN_1095; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1097 = 5'h1f == IFIDrs2 ? Regs_31 : _GEN_1096; // @[cpu.scala 167:{15,15}]
  wire [63:0] _GEN_1099 = bypassBFromWB ? MEMWBValue : _GEN_1097; // @[cpu.scala 163:33 165:11 168:11]
  wire [63:0] _GEN_1101 = bypassBFromMEM ? EXMEMALUOut : _GEN_1099; // @[cpu.scala 160:34 162:11]
  wire [63:0] _GEN_1103 = bypassBFromEX ? _B_T_1 : _GEN_1101; // @[cpu.scala 157:27 159:11]
  wire [63:0] B = ~stall ? _GEN_1103 : 64'h0; // @[cpu.scala 117:27]
  wire  takeBranch = IFIDop == 7'h63 & IFID_funct3 == 3'h0 & A == B; // @[cpu.scala 109:64]
  wire [63:0] _IFIDIR_T = {{2'd0}, PC[63:2]}; // @[cpu.scala 121:31]
  wire [31:0] _GEN_1 = 10'h1 == _IFIDIR_T[9:0] ? IMemory_1 : IMemory_0; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_2 = 10'h2 == _IFIDIR_T[9:0] ? IMemory_2 : _GEN_1; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_3 = 10'h3 == _IFIDIR_T[9:0] ? IMemory_3 : _GEN_2; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_4 = 10'h4 == _IFIDIR_T[9:0] ? IMemory_4 : _GEN_3; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_5 = 10'h5 == _IFIDIR_T[9:0] ? IMemory_5 : _GEN_4; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_6 = 10'h6 == _IFIDIR_T[9:0] ? IMemory_6 : _GEN_5; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_7 = 10'h7 == _IFIDIR_T[9:0] ? IMemory_7 : _GEN_6; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_8 = 10'h8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_7; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_9 = 10'h9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_8; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_10 = 10'ha == _IFIDIR_T[9:0] ? 32'h0 : _GEN_9; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_11 = 10'hb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_10; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_12 = 10'hc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_11; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_13 = 10'hd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_12; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_14 = 10'he == _IFIDIR_T[9:0] ? 32'h0 : _GEN_13; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_15 = 10'hf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_14; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_16 = 10'h10 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_15; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_17 = 10'h11 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_16; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_18 = 10'h12 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_17; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_19 = 10'h13 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_18; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_20 = 10'h14 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_19; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_21 = 10'h15 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_20; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_22 = 10'h16 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_21; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_23 = 10'h17 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_22; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_24 = 10'h18 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_23; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_25 = 10'h19 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_24; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_26 = 10'h1a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_25; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_27 = 10'h1b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_26; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_28 = 10'h1c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_27; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_29 = 10'h1d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_28; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_30 = 10'h1e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_29; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_31 = 10'h1f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_30; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_32 = 10'h20 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_31; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_33 = 10'h21 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_32; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_34 = 10'h22 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_33; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_35 = 10'h23 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_34; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_36 = 10'h24 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_35; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_37 = 10'h25 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_36; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_38 = 10'h26 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_37; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_39 = 10'h27 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_38; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_40 = 10'h28 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_39; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_41 = 10'h29 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_40; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_42 = 10'h2a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_41; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_43 = 10'h2b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_42; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_44 = 10'h2c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_43; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_45 = 10'h2d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_44; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_46 = 10'h2e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_45; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_47 = 10'h2f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_46; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_48 = 10'h30 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_47; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_49 = 10'h31 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_48; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_50 = 10'h32 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_49; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_51 = 10'h33 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_50; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_52 = 10'h34 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_51; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_53 = 10'h35 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_52; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_54 = 10'h36 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_53; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_55 = 10'h37 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_54; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_56 = 10'h38 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_55; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_57 = 10'h39 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_56; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_58 = 10'h3a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_57; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_59 = 10'h3b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_58; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_60 = 10'h3c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_59; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_61 = 10'h3d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_60; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_62 = 10'h3e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_61; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_63 = 10'h3f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_62; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_64 = 10'h40 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_63; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_65 = 10'h41 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_64; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_66 = 10'h42 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_65; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_67 = 10'h43 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_66; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_68 = 10'h44 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_67; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_69 = 10'h45 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_68; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_70 = 10'h46 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_69; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_71 = 10'h47 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_70; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_72 = 10'h48 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_71; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_73 = 10'h49 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_72; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_74 = 10'h4a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_73; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_75 = 10'h4b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_74; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_76 = 10'h4c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_75; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_77 = 10'h4d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_76; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_78 = 10'h4e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_77; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_79 = 10'h4f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_78; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_80 = 10'h50 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_79; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_81 = 10'h51 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_80; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_82 = 10'h52 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_81; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_83 = 10'h53 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_82; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_84 = 10'h54 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_83; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_85 = 10'h55 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_84; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_86 = 10'h56 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_85; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_87 = 10'h57 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_86; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_88 = 10'h58 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_87; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_89 = 10'h59 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_88; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_90 = 10'h5a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_89; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_91 = 10'h5b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_90; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_92 = 10'h5c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_91; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_93 = 10'h5d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_92; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_94 = 10'h5e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_93; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_95 = 10'h5f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_94; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_96 = 10'h60 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_95; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_97 = 10'h61 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_96; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_98 = 10'h62 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_97; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_99 = 10'h63 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_98; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_100 = 10'h64 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_99; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_101 = 10'h65 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_100; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_102 = 10'h66 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_101; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_103 = 10'h67 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_102; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_104 = 10'h68 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_103; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_105 = 10'h69 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_104; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_106 = 10'h6a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_105; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_107 = 10'h6b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_106; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_108 = 10'h6c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_107; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_109 = 10'h6d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_108; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_110 = 10'h6e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_109; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_111 = 10'h6f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_110; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_112 = 10'h70 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_111; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_113 = 10'h71 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_112; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_114 = 10'h72 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_113; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_115 = 10'h73 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_114; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_116 = 10'h74 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_115; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_117 = 10'h75 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_116; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_118 = 10'h76 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_117; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_119 = 10'h77 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_118; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_120 = 10'h78 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_119; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_121 = 10'h79 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_120; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_122 = 10'h7a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_121; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_123 = 10'h7b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_122; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_124 = 10'h7c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_123; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_125 = 10'h7d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_124; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_126 = 10'h7e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_125; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_127 = 10'h7f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_126; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_128 = 10'h80 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_127; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_129 = 10'h81 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_128; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_130 = 10'h82 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_129; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_131 = 10'h83 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_130; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_132 = 10'h84 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_131; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_133 = 10'h85 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_132; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_134 = 10'h86 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_133; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_135 = 10'h87 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_134; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_136 = 10'h88 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_135; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_137 = 10'h89 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_136; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_138 = 10'h8a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_137; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_139 = 10'h8b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_138; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_140 = 10'h8c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_139; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_141 = 10'h8d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_140; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_142 = 10'h8e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_141; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_143 = 10'h8f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_142; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_144 = 10'h90 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_143; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_145 = 10'h91 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_144; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_146 = 10'h92 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_145; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_147 = 10'h93 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_146; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_148 = 10'h94 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_147; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_149 = 10'h95 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_148; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_150 = 10'h96 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_149; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_151 = 10'h97 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_150; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_152 = 10'h98 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_151; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_153 = 10'h99 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_152; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_154 = 10'h9a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_153; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_155 = 10'h9b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_154; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_156 = 10'h9c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_155; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_157 = 10'h9d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_156; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_158 = 10'h9e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_157; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_159 = 10'h9f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_158; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_160 = 10'ha0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_159; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_161 = 10'ha1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_160; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_162 = 10'ha2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_161; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_163 = 10'ha3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_162; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_164 = 10'ha4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_163; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_165 = 10'ha5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_164; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_166 = 10'ha6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_165; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_167 = 10'ha7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_166; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_168 = 10'ha8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_167; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_169 = 10'ha9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_168; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_170 = 10'haa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_169; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_171 = 10'hab == _IFIDIR_T[9:0] ? 32'h0 : _GEN_170; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_172 = 10'hac == _IFIDIR_T[9:0] ? 32'h0 : _GEN_171; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_173 = 10'had == _IFIDIR_T[9:0] ? 32'h0 : _GEN_172; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_174 = 10'hae == _IFIDIR_T[9:0] ? 32'h0 : _GEN_173; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_175 = 10'haf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_174; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_176 = 10'hb0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_175; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_177 = 10'hb1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_176; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_178 = 10'hb2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_177; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_179 = 10'hb3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_178; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_180 = 10'hb4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_179; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_181 = 10'hb5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_180; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_182 = 10'hb6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_181; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_183 = 10'hb7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_182; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_184 = 10'hb8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_183; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_185 = 10'hb9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_184; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_186 = 10'hba == _IFIDIR_T[9:0] ? 32'h0 : _GEN_185; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_187 = 10'hbb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_186; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_188 = 10'hbc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_187; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_189 = 10'hbd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_188; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_190 = 10'hbe == _IFIDIR_T[9:0] ? 32'h0 : _GEN_189; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_191 = 10'hbf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_190; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_192 = 10'hc0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_191; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_193 = 10'hc1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_192; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_194 = 10'hc2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_193; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_195 = 10'hc3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_194; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_196 = 10'hc4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_195; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_197 = 10'hc5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_196; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_198 = 10'hc6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_197; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_199 = 10'hc7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_198; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_200 = 10'hc8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_199; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_201 = 10'hc9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_200; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_202 = 10'hca == _IFIDIR_T[9:0] ? 32'h0 : _GEN_201; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_203 = 10'hcb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_202; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_204 = 10'hcc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_203; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_205 = 10'hcd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_204; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_206 = 10'hce == _IFIDIR_T[9:0] ? 32'h0 : _GEN_205; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_207 = 10'hcf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_206; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_208 = 10'hd0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_207; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_209 = 10'hd1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_208; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_210 = 10'hd2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_209; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_211 = 10'hd3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_210; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_212 = 10'hd4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_211; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_213 = 10'hd5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_212; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_214 = 10'hd6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_213; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_215 = 10'hd7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_214; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_216 = 10'hd8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_215; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_217 = 10'hd9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_216; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_218 = 10'hda == _IFIDIR_T[9:0] ? 32'h0 : _GEN_217; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_219 = 10'hdb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_218; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_220 = 10'hdc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_219; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_221 = 10'hdd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_220; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_222 = 10'hde == _IFIDIR_T[9:0] ? 32'h0 : _GEN_221; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_223 = 10'hdf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_222; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_224 = 10'he0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_223; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_225 = 10'he1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_224; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_226 = 10'he2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_225; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_227 = 10'he3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_226; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_228 = 10'he4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_227; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_229 = 10'he5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_228; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_230 = 10'he6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_229; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_231 = 10'he7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_230; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_232 = 10'he8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_231; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_233 = 10'he9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_232; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_234 = 10'hea == _IFIDIR_T[9:0] ? 32'h0 : _GEN_233; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_235 = 10'heb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_234; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_236 = 10'hec == _IFIDIR_T[9:0] ? 32'h0 : _GEN_235; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_237 = 10'hed == _IFIDIR_T[9:0] ? 32'h0 : _GEN_236; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_238 = 10'hee == _IFIDIR_T[9:0] ? 32'h0 : _GEN_237; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_239 = 10'hef == _IFIDIR_T[9:0] ? 32'h0 : _GEN_238; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_240 = 10'hf0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_239; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_241 = 10'hf1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_240; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_242 = 10'hf2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_241; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_243 = 10'hf3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_242; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_244 = 10'hf4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_243; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_245 = 10'hf5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_244; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_246 = 10'hf6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_245; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_247 = 10'hf7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_246; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_248 = 10'hf8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_247; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_249 = 10'hf9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_248; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_250 = 10'hfa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_249; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_251 = 10'hfb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_250; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_252 = 10'hfc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_251; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_253 = 10'hfd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_252; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_254 = 10'hfe == _IFIDIR_T[9:0] ? 32'h0 : _GEN_253; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_255 = 10'hff == _IFIDIR_T[9:0] ? 32'h0 : _GEN_254; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_256 = 10'h100 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_255; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_257 = 10'h101 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_256; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_258 = 10'h102 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_257; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_259 = 10'h103 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_258; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_260 = 10'h104 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_259; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_261 = 10'h105 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_260; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_262 = 10'h106 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_261; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_263 = 10'h107 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_262; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_264 = 10'h108 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_263; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_265 = 10'h109 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_264; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_266 = 10'h10a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_265; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_267 = 10'h10b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_266; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_268 = 10'h10c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_267; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_269 = 10'h10d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_268; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_270 = 10'h10e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_269; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_271 = 10'h10f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_270; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_272 = 10'h110 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_271; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_273 = 10'h111 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_272; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_274 = 10'h112 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_273; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_275 = 10'h113 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_274; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_276 = 10'h114 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_275; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_277 = 10'h115 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_276; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_278 = 10'h116 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_277; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_279 = 10'h117 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_278; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_280 = 10'h118 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_279; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_281 = 10'h119 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_280; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_282 = 10'h11a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_281; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_283 = 10'h11b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_282; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_284 = 10'h11c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_283; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_285 = 10'h11d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_284; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_286 = 10'h11e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_285; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_287 = 10'h11f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_286; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_288 = 10'h120 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_287; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_289 = 10'h121 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_288; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_290 = 10'h122 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_289; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_291 = 10'h123 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_290; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_292 = 10'h124 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_291; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_293 = 10'h125 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_292; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_294 = 10'h126 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_293; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_295 = 10'h127 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_294; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_296 = 10'h128 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_295; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_297 = 10'h129 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_296; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_298 = 10'h12a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_297; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_299 = 10'h12b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_298; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_300 = 10'h12c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_299; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_301 = 10'h12d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_300; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_302 = 10'h12e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_301; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_303 = 10'h12f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_302; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_304 = 10'h130 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_303; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_305 = 10'h131 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_304; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_306 = 10'h132 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_305; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_307 = 10'h133 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_306; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_308 = 10'h134 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_307; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_309 = 10'h135 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_308; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_310 = 10'h136 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_309; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_311 = 10'h137 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_310; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_312 = 10'h138 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_311; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_313 = 10'h139 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_312; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_314 = 10'h13a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_313; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_315 = 10'h13b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_314; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_316 = 10'h13c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_315; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_317 = 10'h13d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_316; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_318 = 10'h13e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_317; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_319 = 10'h13f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_318; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_320 = 10'h140 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_319; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_321 = 10'h141 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_320; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_322 = 10'h142 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_321; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_323 = 10'h143 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_322; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_324 = 10'h144 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_323; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_325 = 10'h145 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_324; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_326 = 10'h146 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_325; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_327 = 10'h147 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_326; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_328 = 10'h148 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_327; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_329 = 10'h149 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_328; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_330 = 10'h14a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_329; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_331 = 10'h14b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_330; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_332 = 10'h14c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_331; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_333 = 10'h14d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_332; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_334 = 10'h14e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_333; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_335 = 10'h14f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_334; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_336 = 10'h150 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_335; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_337 = 10'h151 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_336; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_338 = 10'h152 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_337; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_339 = 10'h153 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_338; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_340 = 10'h154 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_339; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_341 = 10'h155 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_340; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_342 = 10'h156 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_341; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_343 = 10'h157 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_342; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_344 = 10'h158 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_343; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_345 = 10'h159 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_344; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_346 = 10'h15a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_345; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_347 = 10'h15b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_346; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_348 = 10'h15c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_347; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_349 = 10'h15d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_348; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_350 = 10'h15e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_349; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_351 = 10'h15f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_350; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_352 = 10'h160 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_351; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_353 = 10'h161 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_352; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_354 = 10'h162 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_353; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_355 = 10'h163 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_354; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_356 = 10'h164 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_355; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_357 = 10'h165 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_356; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_358 = 10'h166 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_357; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_359 = 10'h167 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_358; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_360 = 10'h168 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_359; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_361 = 10'h169 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_360; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_362 = 10'h16a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_361; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_363 = 10'h16b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_362; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_364 = 10'h16c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_363; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_365 = 10'h16d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_364; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_366 = 10'h16e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_365; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_367 = 10'h16f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_366; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_368 = 10'h170 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_367; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_369 = 10'h171 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_368; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_370 = 10'h172 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_369; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_371 = 10'h173 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_370; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_372 = 10'h174 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_371; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_373 = 10'h175 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_372; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_374 = 10'h176 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_373; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_375 = 10'h177 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_374; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_376 = 10'h178 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_375; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_377 = 10'h179 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_376; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_378 = 10'h17a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_377; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_379 = 10'h17b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_378; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_380 = 10'h17c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_379; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_381 = 10'h17d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_380; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_382 = 10'h17e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_381; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_383 = 10'h17f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_382; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_384 = 10'h180 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_383; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_385 = 10'h181 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_384; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_386 = 10'h182 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_385; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_387 = 10'h183 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_386; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_388 = 10'h184 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_387; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_389 = 10'h185 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_388; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_390 = 10'h186 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_389; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_391 = 10'h187 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_390; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_392 = 10'h188 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_391; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_393 = 10'h189 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_392; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_394 = 10'h18a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_393; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_395 = 10'h18b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_394; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_396 = 10'h18c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_395; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_397 = 10'h18d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_396; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_398 = 10'h18e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_397; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_399 = 10'h18f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_398; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_400 = 10'h190 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_399; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_401 = 10'h191 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_400; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_402 = 10'h192 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_401; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_403 = 10'h193 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_402; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_404 = 10'h194 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_403; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_405 = 10'h195 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_404; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_406 = 10'h196 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_405; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_407 = 10'h197 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_406; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_408 = 10'h198 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_407; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_409 = 10'h199 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_408; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_410 = 10'h19a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_409; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_411 = 10'h19b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_410; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_412 = 10'h19c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_411; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_413 = 10'h19d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_412; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_414 = 10'h19e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_413; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_415 = 10'h19f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_414; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_416 = 10'h1a0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_415; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_417 = 10'h1a1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_416; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_418 = 10'h1a2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_417; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_419 = 10'h1a3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_418; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_420 = 10'h1a4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_419; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_421 = 10'h1a5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_420; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_422 = 10'h1a6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_421; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_423 = 10'h1a7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_422; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_424 = 10'h1a8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_423; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_425 = 10'h1a9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_424; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_426 = 10'h1aa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_425; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_427 = 10'h1ab == _IFIDIR_T[9:0] ? 32'h0 : _GEN_426; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_428 = 10'h1ac == _IFIDIR_T[9:0] ? 32'h0 : _GEN_427; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_429 = 10'h1ad == _IFIDIR_T[9:0] ? 32'h0 : _GEN_428; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_430 = 10'h1ae == _IFIDIR_T[9:0] ? 32'h0 : _GEN_429; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_431 = 10'h1af == _IFIDIR_T[9:0] ? 32'h0 : _GEN_430; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_432 = 10'h1b0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_431; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_433 = 10'h1b1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_432; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_434 = 10'h1b2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_433; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_435 = 10'h1b3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_434; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_436 = 10'h1b4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_435; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_437 = 10'h1b5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_436; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_438 = 10'h1b6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_437; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_439 = 10'h1b7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_438; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_440 = 10'h1b8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_439; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_441 = 10'h1b9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_440; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_442 = 10'h1ba == _IFIDIR_T[9:0] ? 32'h0 : _GEN_441; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_443 = 10'h1bb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_442; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_444 = 10'h1bc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_443; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_445 = 10'h1bd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_444; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_446 = 10'h1be == _IFIDIR_T[9:0] ? 32'h0 : _GEN_445; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_447 = 10'h1bf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_446; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_448 = 10'h1c0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_447; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_449 = 10'h1c1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_448; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_450 = 10'h1c2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_449; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_451 = 10'h1c3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_450; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_452 = 10'h1c4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_451; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_453 = 10'h1c5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_452; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_454 = 10'h1c6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_453; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_455 = 10'h1c7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_454; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_456 = 10'h1c8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_455; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_457 = 10'h1c9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_456; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_458 = 10'h1ca == _IFIDIR_T[9:0] ? 32'h0 : _GEN_457; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_459 = 10'h1cb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_458; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_460 = 10'h1cc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_459; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_461 = 10'h1cd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_460; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_462 = 10'h1ce == _IFIDIR_T[9:0] ? 32'h0 : _GEN_461; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_463 = 10'h1cf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_462; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_464 = 10'h1d0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_463; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_465 = 10'h1d1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_464; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_466 = 10'h1d2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_465; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_467 = 10'h1d3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_466; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_468 = 10'h1d4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_467; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_469 = 10'h1d5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_468; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_470 = 10'h1d6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_469; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_471 = 10'h1d7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_470; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_472 = 10'h1d8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_471; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_473 = 10'h1d9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_472; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_474 = 10'h1da == _IFIDIR_T[9:0] ? 32'h0 : _GEN_473; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_475 = 10'h1db == _IFIDIR_T[9:0] ? 32'h0 : _GEN_474; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_476 = 10'h1dc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_475; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_477 = 10'h1dd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_476; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_478 = 10'h1de == _IFIDIR_T[9:0] ? 32'h0 : _GEN_477; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_479 = 10'h1df == _IFIDIR_T[9:0] ? 32'h0 : _GEN_478; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_480 = 10'h1e0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_479; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_481 = 10'h1e1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_480; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_482 = 10'h1e2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_481; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_483 = 10'h1e3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_482; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_484 = 10'h1e4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_483; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_485 = 10'h1e5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_484; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_486 = 10'h1e6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_485; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_487 = 10'h1e7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_486; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_488 = 10'h1e8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_487; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_489 = 10'h1e9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_488; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_490 = 10'h1ea == _IFIDIR_T[9:0] ? 32'h0 : _GEN_489; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_491 = 10'h1eb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_490; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_492 = 10'h1ec == _IFIDIR_T[9:0] ? 32'h0 : _GEN_491; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_493 = 10'h1ed == _IFIDIR_T[9:0] ? 32'h0 : _GEN_492; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_494 = 10'h1ee == _IFIDIR_T[9:0] ? 32'h0 : _GEN_493; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_495 = 10'h1ef == _IFIDIR_T[9:0] ? 32'h0 : _GEN_494; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_496 = 10'h1f0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_495; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_497 = 10'h1f1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_496; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_498 = 10'h1f2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_497; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_499 = 10'h1f3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_498; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_500 = 10'h1f4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_499; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_501 = 10'h1f5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_500; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_502 = 10'h1f6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_501; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_503 = 10'h1f7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_502; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_504 = 10'h1f8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_503; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_505 = 10'h1f9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_504; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_506 = 10'h1fa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_505; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_507 = 10'h1fb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_506; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_508 = 10'h1fc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_507; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_509 = 10'h1fd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_508; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_510 = 10'h1fe == _IFIDIR_T[9:0] ? 32'h0 : _GEN_509; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_511 = 10'h1ff == _IFIDIR_T[9:0] ? 32'h0 : _GEN_510; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_512 = 10'h200 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_511; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_513 = 10'h201 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_512; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_514 = 10'h202 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_513; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_515 = 10'h203 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_514; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_516 = 10'h204 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_515; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_517 = 10'h205 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_516; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_518 = 10'h206 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_517; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_519 = 10'h207 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_518; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_520 = 10'h208 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_519; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_521 = 10'h209 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_520; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_522 = 10'h20a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_521; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_523 = 10'h20b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_522; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_524 = 10'h20c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_523; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_525 = 10'h20d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_524; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_526 = 10'h20e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_525; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_527 = 10'h20f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_526; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_528 = 10'h210 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_527; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_529 = 10'h211 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_528; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_530 = 10'h212 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_529; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_531 = 10'h213 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_530; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_532 = 10'h214 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_531; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_533 = 10'h215 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_532; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_534 = 10'h216 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_533; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_535 = 10'h217 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_534; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_536 = 10'h218 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_535; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_537 = 10'h219 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_536; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_538 = 10'h21a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_537; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_539 = 10'h21b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_538; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_540 = 10'h21c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_539; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_541 = 10'h21d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_540; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_542 = 10'h21e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_541; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_543 = 10'h21f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_542; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_544 = 10'h220 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_543; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_545 = 10'h221 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_544; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_546 = 10'h222 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_545; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_547 = 10'h223 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_546; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_548 = 10'h224 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_547; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_549 = 10'h225 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_548; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_550 = 10'h226 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_549; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_551 = 10'h227 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_550; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_552 = 10'h228 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_551; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_553 = 10'h229 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_552; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_554 = 10'h22a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_553; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_555 = 10'h22b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_554; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_556 = 10'h22c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_555; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_557 = 10'h22d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_556; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_558 = 10'h22e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_557; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_559 = 10'h22f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_558; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_560 = 10'h230 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_559; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_561 = 10'h231 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_560; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_562 = 10'h232 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_561; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_563 = 10'h233 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_562; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_564 = 10'h234 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_563; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_565 = 10'h235 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_564; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_566 = 10'h236 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_565; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_567 = 10'h237 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_566; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_568 = 10'h238 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_567; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_569 = 10'h239 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_568; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_570 = 10'h23a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_569; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_571 = 10'h23b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_570; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_572 = 10'h23c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_571; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_573 = 10'h23d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_572; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_574 = 10'h23e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_573; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_575 = 10'h23f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_574; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_576 = 10'h240 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_575; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_577 = 10'h241 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_576; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_578 = 10'h242 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_577; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_579 = 10'h243 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_578; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_580 = 10'h244 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_579; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_581 = 10'h245 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_580; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_582 = 10'h246 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_581; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_583 = 10'h247 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_582; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_584 = 10'h248 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_583; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_585 = 10'h249 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_584; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_586 = 10'h24a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_585; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_587 = 10'h24b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_586; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_588 = 10'h24c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_587; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_589 = 10'h24d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_588; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_590 = 10'h24e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_589; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_591 = 10'h24f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_590; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_592 = 10'h250 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_591; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_593 = 10'h251 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_592; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_594 = 10'h252 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_593; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_595 = 10'h253 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_594; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_596 = 10'h254 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_595; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_597 = 10'h255 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_596; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_598 = 10'h256 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_597; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_599 = 10'h257 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_598; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_600 = 10'h258 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_599; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_601 = 10'h259 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_600; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_602 = 10'h25a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_601; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_603 = 10'h25b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_602; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_604 = 10'h25c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_603; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_605 = 10'h25d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_604; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_606 = 10'h25e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_605; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_607 = 10'h25f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_606; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_608 = 10'h260 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_607; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_609 = 10'h261 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_608; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_610 = 10'h262 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_609; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_611 = 10'h263 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_610; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_612 = 10'h264 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_611; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_613 = 10'h265 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_612; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_614 = 10'h266 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_613; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_615 = 10'h267 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_614; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_616 = 10'h268 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_615; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_617 = 10'h269 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_616; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_618 = 10'h26a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_617; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_619 = 10'h26b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_618; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_620 = 10'h26c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_619; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_621 = 10'h26d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_620; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_622 = 10'h26e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_621; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_623 = 10'h26f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_622; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_624 = 10'h270 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_623; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_625 = 10'h271 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_624; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_626 = 10'h272 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_625; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_627 = 10'h273 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_626; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_628 = 10'h274 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_627; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_629 = 10'h275 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_628; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_630 = 10'h276 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_629; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_631 = 10'h277 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_630; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_632 = 10'h278 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_631; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_633 = 10'h279 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_632; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_634 = 10'h27a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_633; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_635 = 10'h27b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_634; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_636 = 10'h27c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_635; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_637 = 10'h27d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_636; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_638 = 10'h27e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_637; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_639 = 10'h27f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_638; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_640 = 10'h280 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_639; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_641 = 10'h281 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_640; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_642 = 10'h282 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_641; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_643 = 10'h283 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_642; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_644 = 10'h284 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_643; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_645 = 10'h285 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_644; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_646 = 10'h286 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_645; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_647 = 10'h287 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_646; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_648 = 10'h288 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_647; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_649 = 10'h289 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_648; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_650 = 10'h28a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_649; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_651 = 10'h28b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_650; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_652 = 10'h28c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_651; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_653 = 10'h28d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_652; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_654 = 10'h28e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_653; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_655 = 10'h28f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_654; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_656 = 10'h290 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_655; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_657 = 10'h291 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_656; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_658 = 10'h292 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_657; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_659 = 10'h293 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_658; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_660 = 10'h294 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_659; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_661 = 10'h295 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_660; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_662 = 10'h296 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_661; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_663 = 10'h297 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_662; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_664 = 10'h298 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_663; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_665 = 10'h299 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_664; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_666 = 10'h29a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_665; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_667 = 10'h29b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_666; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_668 = 10'h29c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_667; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_669 = 10'h29d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_668; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_670 = 10'h29e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_669; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_671 = 10'h29f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_670; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_672 = 10'h2a0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_671; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_673 = 10'h2a1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_672; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_674 = 10'h2a2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_673; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_675 = 10'h2a3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_674; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_676 = 10'h2a4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_675; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_677 = 10'h2a5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_676; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_678 = 10'h2a6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_677; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_679 = 10'h2a7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_678; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_680 = 10'h2a8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_679; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_681 = 10'h2a9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_680; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_682 = 10'h2aa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_681; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_683 = 10'h2ab == _IFIDIR_T[9:0] ? 32'h0 : _GEN_682; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_684 = 10'h2ac == _IFIDIR_T[9:0] ? 32'h0 : _GEN_683; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_685 = 10'h2ad == _IFIDIR_T[9:0] ? 32'h0 : _GEN_684; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_686 = 10'h2ae == _IFIDIR_T[9:0] ? 32'h0 : _GEN_685; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_687 = 10'h2af == _IFIDIR_T[9:0] ? 32'h0 : _GEN_686; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_688 = 10'h2b0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_687; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_689 = 10'h2b1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_688; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_690 = 10'h2b2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_689; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_691 = 10'h2b3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_690; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_692 = 10'h2b4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_691; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_693 = 10'h2b5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_692; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_694 = 10'h2b6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_693; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_695 = 10'h2b7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_694; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_696 = 10'h2b8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_695; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_697 = 10'h2b9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_696; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_698 = 10'h2ba == _IFIDIR_T[9:0] ? 32'h0 : _GEN_697; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_699 = 10'h2bb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_698; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_700 = 10'h2bc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_699; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_701 = 10'h2bd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_700; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_702 = 10'h2be == _IFIDIR_T[9:0] ? 32'h0 : _GEN_701; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_703 = 10'h2bf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_702; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_704 = 10'h2c0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_703; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_705 = 10'h2c1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_704; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_706 = 10'h2c2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_705; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_707 = 10'h2c3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_706; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_708 = 10'h2c4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_707; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_709 = 10'h2c5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_708; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_710 = 10'h2c6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_709; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_711 = 10'h2c7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_710; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_712 = 10'h2c8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_711; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_713 = 10'h2c9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_712; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_714 = 10'h2ca == _IFIDIR_T[9:0] ? 32'h0 : _GEN_713; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_715 = 10'h2cb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_714; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_716 = 10'h2cc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_715; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_717 = 10'h2cd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_716; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_718 = 10'h2ce == _IFIDIR_T[9:0] ? 32'h0 : _GEN_717; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_719 = 10'h2cf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_718; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_720 = 10'h2d0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_719; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_721 = 10'h2d1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_720; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_722 = 10'h2d2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_721; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_723 = 10'h2d3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_722; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_724 = 10'h2d4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_723; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_725 = 10'h2d5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_724; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_726 = 10'h2d6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_725; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_727 = 10'h2d7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_726; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_728 = 10'h2d8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_727; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_729 = 10'h2d9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_728; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_730 = 10'h2da == _IFIDIR_T[9:0] ? 32'h0 : _GEN_729; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_731 = 10'h2db == _IFIDIR_T[9:0] ? 32'h0 : _GEN_730; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_732 = 10'h2dc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_731; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_733 = 10'h2dd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_732; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_734 = 10'h2de == _IFIDIR_T[9:0] ? 32'h0 : _GEN_733; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_735 = 10'h2df == _IFIDIR_T[9:0] ? 32'h0 : _GEN_734; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_736 = 10'h2e0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_735; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_737 = 10'h2e1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_736; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_738 = 10'h2e2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_737; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_739 = 10'h2e3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_738; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_740 = 10'h2e4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_739; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_741 = 10'h2e5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_740; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_742 = 10'h2e6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_741; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_743 = 10'h2e7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_742; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_744 = 10'h2e8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_743; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_745 = 10'h2e9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_744; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_746 = 10'h2ea == _IFIDIR_T[9:0] ? 32'h0 : _GEN_745; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_747 = 10'h2eb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_746; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_748 = 10'h2ec == _IFIDIR_T[9:0] ? 32'h0 : _GEN_747; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_749 = 10'h2ed == _IFIDIR_T[9:0] ? 32'h0 : _GEN_748; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_750 = 10'h2ee == _IFIDIR_T[9:0] ? 32'h0 : _GEN_749; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_751 = 10'h2ef == _IFIDIR_T[9:0] ? 32'h0 : _GEN_750; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_752 = 10'h2f0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_751; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_753 = 10'h2f1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_752; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_754 = 10'h2f2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_753; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_755 = 10'h2f3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_754; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_756 = 10'h2f4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_755; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_757 = 10'h2f5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_756; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_758 = 10'h2f6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_757; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_759 = 10'h2f7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_758; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_760 = 10'h2f8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_759; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_761 = 10'h2f9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_760; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_762 = 10'h2fa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_761; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_763 = 10'h2fb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_762; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_764 = 10'h2fc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_763; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_765 = 10'h2fd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_764; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_766 = 10'h2fe == _IFIDIR_T[9:0] ? 32'h0 : _GEN_765; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_767 = 10'h2ff == _IFIDIR_T[9:0] ? 32'h0 : _GEN_766; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_768 = 10'h300 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_767; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_769 = 10'h301 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_768; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_770 = 10'h302 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_769; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_771 = 10'h303 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_770; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_772 = 10'h304 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_771; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_773 = 10'h305 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_772; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_774 = 10'h306 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_773; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_775 = 10'h307 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_774; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_776 = 10'h308 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_775; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_777 = 10'h309 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_776; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_778 = 10'h30a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_777; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_779 = 10'h30b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_778; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_780 = 10'h30c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_779; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_781 = 10'h30d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_780; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_782 = 10'h30e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_781; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_783 = 10'h30f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_782; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_784 = 10'h310 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_783; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_785 = 10'h311 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_784; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_786 = 10'h312 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_785; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_787 = 10'h313 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_786; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_788 = 10'h314 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_787; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_789 = 10'h315 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_788; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_790 = 10'h316 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_789; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_791 = 10'h317 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_790; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_792 = 10'h318 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_791; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_793 = 10'h319 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_792; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_794 = 10'h31a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_793; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_795 = 10'h31b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_794; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_796 = 10'h31c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_795; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_797 = 10'h31d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_796; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_798 = 10'h31e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_797; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_799 = 10'h31f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_798; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_800 = 10'h320 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_799; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_801 = 10'h321 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_800; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_802 = 10'h322 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_801; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_803 = 10'h323 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_802; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_804 = 10'h324 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_803; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_805 = 10'h325 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_804; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_806 = 10'h326 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_805; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_807 = 10'h327 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_806; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_808 = 10'h328 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_807; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_809 = 10'h329 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_808; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_810 = 10'h32a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_809; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_811 = 10'h32b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_810; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_812 = 10'h32c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_811; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_813 = 10'h32d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_812; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_814 = 10'h32e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_813; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_815 = 10'h32f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_814; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_816 = 10'h330 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_815; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_817 = 10'h331 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_816; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_818 = 10'h332 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_817; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_819 = 10'h333 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_818; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_820 = 10'h334 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_819; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_821 = 10'h335 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_820; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_822 = 10'h336 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_821; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_823 = 10'h337 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_822; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_824 = 10'h338 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_823; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_825 = 10'h339 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_824; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_826 = 10'h33a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_825; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_827 = 10'h33b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_826; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_828 = 10'h33c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_827; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_829 = 10'h33d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_828; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_830 = 10'h33e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_829; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_831 = 10'h33f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_830; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_832 = 10'h340 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_831; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_833 = 10'h341 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_832; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_834 = 10'h342 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_833; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_835 = 10'h343 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_834; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_836 = 10'h344 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_835; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_837 = 10'h345 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_836; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_838 = 10'h346 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_837; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_839 = 10'h347 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_838; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_840 = 10'h348 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_839; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_841 = 10'h349 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_840; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_842 = 10'h34a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_841; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_843 = 10'h34b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_842; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_844 = 10'h34c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_843; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_845 = 10'h34d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_844; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_846 = 10'h34e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_845; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_847 = 10'h34f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_846; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_848 = 10'h350 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_847; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_849 = 10'h351 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_848; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_850 = 10'h352 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_849; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_851 = 10'h353 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_850; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_852 = 10'h354 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_851; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_853 = 10'h355 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_852; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_854 = 10'h356 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_853; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_855 = 10'h357 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_854; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_856 = 10'h358 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_855; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_857 = 10'h359 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_856; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_858 = 10'h35a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_857; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_859 = 10'h35b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_858; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_860 = 10'h35c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_859; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_861 = 10'h35d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_860; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_862 = 10'h35e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_861; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_863 = 10'h35f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_862; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_864 = 10'h360 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_863; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_865 = 10'h361 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_864; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_866 = 10'h362 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_865; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_867 = 10'h363 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_866; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_868 = 10'h364 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_867; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_869 = 10'h365 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_868; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_870 = 10'h366 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_869; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_871 = 10'h367 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_870; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_872 = 10'h368 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_871; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_873 = 10'h369 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_872; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_874 = 10'h36a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_873; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_875 = 10'h36b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_874; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_876 = 10'h36c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_875; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_877 = 10'h36d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_876; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_878 = 10'h36e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_877; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_879 = 10'h36f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_878; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_880 = 10'h370 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_879; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_881 = 10'h371 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_880; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_882 = 10'h372 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_881; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_883 = 10'h373 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_882; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_884 = 10'h374 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_883; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_885 = 10'h375 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_884; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_886 = 10'h376 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_885; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_887 = 10'h377 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_886; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_888 = 10'h378 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_887; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_889 = 10'h379 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_888; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_890 = 10'h37a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_889; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_891 = 10'h37b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_890; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_892 = 10'h37c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_891; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_893 = 10'h37d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_892; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_894 = 10'h37e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_893; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_895 = 10'h37f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_894; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_896 = 10'h380 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_895; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_897 = 10'h381 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_896; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_898 = 10'h382 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_897; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_899 = 10'h383 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_898; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_900 = 10'h384 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_899; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_901 = 10'h385 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_900; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_902 = 10'h386 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_901; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_903 = 10'h387 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_902; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_904 = 10'h388 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_903; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_905 = 10'h389 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_904; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_906 = 10'h38a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_905; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_907 = 10'h38b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_906; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_908 = 10'h38c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_907; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_909 = 10'h38d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_908; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_910 = 10'h38e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_909; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_911 = 10'h38f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_910; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_912 = 10'h390 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_911; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_913 = 10'h391 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_912; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_914 = 10'h392 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_913; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_915 = 10'h393 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_914; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_916 = 10'h394 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_915; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_917 = 10'h395 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_916; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_918 = 10'h396 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_917; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_919 = 10'h397 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_918; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_920 = 10'h398 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_919; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_921 = 10'h399 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_920; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_922 = 10'h39a == _IFIDIR_T[9:0] ? 32'h0 : _GEN_921; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_923 = 10'h39b == _IFIDIR_T[9:0] ? 32'h0 : _GEN_922; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_924 = 10'h39c == _IFIDIR_T[9:0] ? 32'h0 : _GEN_923; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_925 = 10'h39d == _IFIDIR_T[9:0] ? 32'h0 : _GEN_924; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_926 = 10'h39e == _IFIDIR_T[9:0] ? 32'h0 : _GEN_925; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_927 = 10'h39f == _IFIDIR_T[9:0] ? 32'h0 : _GEN_926; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_928 = 10'h3a0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_927; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_929 = 10'h3a1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_928; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_930 = 10'h3a2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_929; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_931 = 10'h3a3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_930; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_932 = 10'h3a4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_931; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_933 = 10'h3a5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_932; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_934 = 10'h3a6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_933; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_935 = 10'h3a7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_934; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_936 = 10'h3a8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_935; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_937 = 10'h3a9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_936; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_938 = 10'h3aa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_937; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_939 = 10'h3ab == _IFIDIR_T[9:0] ? 32'h0 : _GEN_938; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_940 = 10'h3ac == _IFIDIR_T[9:0] ? 32'h0 : _GEN_939; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_941 = 10'h3ad == _IFIDIR_T[9:0] ? 32'h0 : _GEN_940; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_942 = 10'h3ae == _IFIDIR_T[9:0] ? 32'h0 : _GEN_941; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_943 = 10'h3af == _IFIDIR_T[9:0] ? 32'h0 : _GEN_942; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_944 = 10'h3b0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_943; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_945 = 10'h3b1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_944; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_946 = 10'h3b2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_945; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_947 = 10'h3b3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_946; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_948 = 10'h3b4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_947; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_949 = 10'h3b5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_948; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_950 = 10'h3b6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_949; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_951 = 10'h3b7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_950; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_952 = 10'h3b8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_951; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_953 = 10'h3b9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_952; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_954 = 10'h3ba == _IFIDIR_T[9:0] ? 32'h0 : _GEN_953; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_955 = 10'h3bb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_954; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_956 = 10'h3bc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_955; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_957 = 10'h3bd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_956; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_958 = 10'h3be == _IFIDIR_T[9:0] ? 32'h0 : _GEN_957; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_959 = 10'h3bf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_958; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_960 = 10'h3c0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_959; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_961 = 10'h3c1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_960; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_962 = 10'h3c2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_961; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_963 = 10'h3c3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_962; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_964 = 10'h3c4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_963; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_965 = 10'h3c5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_964; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_966 = 10'h3c6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_965; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_967 = 10'h3c7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_966; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_968 = 10'h3c8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_967; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_969 = 10'h3c9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_968; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_970 = 10'h3ca == _IFIDIR_T[9:0] ? 32'h0 : _GEN_969; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_971 = 10'h3cb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_970; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_972 = 10'h3cc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_971; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_973 = 10'h3cd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_972; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_974 = 10'h3ce == _IFIDIR_T[9:0] ? 32'h0 : _GEN_973; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_975 = 10'h3cf == _IFIDIR_T[9:0] ? 32'h0 : _GEN_974; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_976 = 10'h3d0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_975; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_977 = 10'h3d1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_976; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_978 = 10'h3d2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_977; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_979 = 10'h3d3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_978; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_980 = 10'h3d4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_979; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_981 = 10'h3d5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_980; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_982 = 10'h3d6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_981; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_983 = 10'h3d7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_982; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_984 = 10'h3d8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_983; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_985 = 10'h3d9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_984; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_986 = 10'h3da == _IFIDIR_T[9:0] ? 32'h0 : _GEN_985; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_987 = 10'h3db == _IFIDIR_T[9:0] ? 32'h0 : _GEN_986; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_988 = 10'h3dc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_987; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_989 = 10'h3dd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_988; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_990 = 10'h3de == _IFIDIR_T[9:0] ? 32'h0 : _GEN_989; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_991 = 10'h3df == _IFIDIR_T[9:0] ? 32'h0 : _GEN_990; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_992 = 10'h3e0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_991; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_993 = 10'h3e1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_992; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_994 = 10'h3e2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_993; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_995 = 10'h3e3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_994; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_996 = 10'h3e4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_995; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_997 = 10'h3e5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_996; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_998 = 10'h3e6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_997; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_999 = 10'h3e7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_998; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1000 = 10'h3e8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_999; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1001 = 10'h3e9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1000; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1002 = 10'h3ea == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1001; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1003 = 10'h3eb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1002; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1004 = 10'h3ec == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1003; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1005 = 10'h3ed == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1004; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1006 = 10'h3ee == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1005; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1007 = 10'h3ef == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1006; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1008 = 10'h3f0 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1007; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1009 = 10'h3f1 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1008; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1010 = 10'h3f2 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1009; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1011 = 10'h3f3 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1010; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1012 = 10'h3f4 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1011; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1013 = 10'h3f5 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1012; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1014 = 10'h3f6 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1013; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1015 = 10'h3f7 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1014; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1016 = 10'h3f8 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1015; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1017 = 10'h3f9 == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1016; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1018 = 10'h3fa == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1017; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1019 = 10'h3fb == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1018; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1020 = 10'h3fc == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1019; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1021 = 10'h3fd == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1020; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1022 = 10'h3fe == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1021; // @[cpu.scala 121:{16,16}]
  wire [31:0] _GEN_1023 = 10'h3ff == _IFIDIR_T[9:0] ? 32'h0 : _GEN_1022; // @[cpu.scala 121:{16,16}]
  wire [63:0] _PC_T_1 = PC + 64'h4; // @[cpu.scala 122:18]
  wire [12:0] _branchTarget_T_5 = {IFIDIR[31],1'h0,IFIDIR[30:25],IFIDIR[11:7]}; // @[cpu.scala 131:11]
  wire [63:0] _GEN_7388 = {{51{_branchTarget_T_5[12]}},_branchTarget_T_5}; // @[cpu.scala 126:42]
  wire [63:0] branchTarget = $signed(CurPC) + $signed(_GEN_7388); // @[cpu.scala 131:19]
  wire [11:0] _EXMEMALUOut_T_2 = IDEXIR[31:20]; // @[cpu.scala 179:53]
  wire [63:0] _GEN_7389 = {{52{_EXMEMALUOut_T_2[11]}},_EXMEMALUOut_T_2}; // @[cpu.scala 179:36]
  wire [63:0] _EXMEMALUOut_T_6 = $signed(IDEXA) + $signed(_GEN_7389); // @[cpu.scala 179:61]
  wire [11:0] _EXMEMALUOut_T_11 = {IDEXIR[31:25],IDEXrd}; // @[cpu.scala 184:9]
  wire [63:0] _GEN_7390 = {{52{_EXMEMALUOut_T_11[11]}},_EXMEMALUOut_T_11}; // @[cpu.scala 181:36]
  wire [63:0] _EXMEMALUOut_T_15 = $signed(IDEXA) + $signed(_GEN_7390); // @[cpu.scala 184:17]
  wire [31:0] _GEN_1118 = 10'h1 == EXMEMALUOut[9:0] ? DMemory_1 : DMemory_0; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1119 = 10'h2 == EXMEMALUOut[9:0] ? DMemory_2 : _GEN_1118; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1120 = 10'h3 == EXMEMALUOut[9:0] ? DMemory_3 : _GEN_1119; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1121 = 10'h4 == EXMEMALUOut[9:0] ? DMemory_4 : _GEN_1120; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1122 = 10'h5 == EXMEMALUOut[9:0] ? DMemory_5 : _GEN_1121; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1123 = 10'h6 == EXMEMALUOut[9:0] ? DMemory_6 : _GEN_1122; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1124 = 10'h7 == EXMEMALUOut[9:0] ? DMemory_7 : _GEN_1123; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1125 = 10'h8 == EXMEMALUOut[9:0] ? DMemory_8 : _GEN_1124; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1126 = 10'h9 == EXMEMALUOut[9:0] ? DMemory_9 : _GEN_1125; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1127 = 10'ha == EXMEMALUOut[9:0] ? DMemory_10 : _GEN_1126; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1128 = 10'hb == EXMEMALUOut[9:0] ? DMemory_11 : _GEN_1127; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1129 = 10'hc == EXMEMALUOut[9:0] ? DMemory_12 : _GEN_1128; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1130 = 10'hd == EXMEMALUOut[9:0] ? DMemory_13 : _GEN_1129; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1131 = 10'he == EXMEMALUOut[9:0] ? DMemory_14 : _GEN_1130; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1132 = 10'hf == EXMEMALUOut[9:0] ? DMemory_15 : _GEN_1131; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1133 = 10'h10 == EXMEMALUOut[9:0] ? DMemory_16 : _GEN_1132; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1134 = 10'h11 == EXMEMALUOut[9:0] ? DMemory_17 : _GEN_1133; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1135 = 10'h12 == EXMEMALUOut[9:0] ? DMemory_18 : _GEN_1134; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1136 = 10'h13 == EXMEMALUOut[9:0] ? DMemory_19 : _GEN_1135; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1137 = 10'h14 == EXMEMALUOut[9:0] ? DMemory_20 : _GEN_1136; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1138 = 10'h15 == EXMEMALUOut[9:0] ? DMemory_21 : _GEN_1137; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1139 = 10'h16 == EXMEMALUOut[9:0] ? DMemory_22 : _GEN_1138; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1140 = 10'h17 == EXMEMALUOut[9:0] ? DMemory_23 : _GEN_1139; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1141 = 10'h18 == EXMEMALUOut[9:0] ? DMemory_24 : _GEN_1140; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1142 = 10'h19 == EXMEMALUOut[9:0] ? DMemory_25 : _GEN_1141; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1143 = 10'h1a == EXMEMALUOut[9:0] ? DMemory_26 : _GEN_1142; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1144 = 10'h1b == EXMEMALUOut[9:0] ? DMemory_27 : _GEN_1143; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1145 = 10'h1c == EXMEMALUOut[9:0] ? DMemory_28 : _GEN_1144; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1146 = 10'h1d == EXMEMALUOut[9:0] ? DMemory_29 : _GEN_1145; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1147 = 10'h1e == EXMEMALUOut[9:0] ? DMemory_30 : _GEN_1146; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1148 = 10'h1f == EXMEMALUOut[9:0] ? DMemory_31 : _GEN_1147; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1149 = 10'h20 == EXMEMALUOut[9:0] ? DMemory_32 : _GEN_1148; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1150 = 10'h21 == EXMEMALUOut[9:0] ? DMemory_33 : _GEN_1149; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1151 = 10'h22 == EXMEMALUOut[9:0] ? DMemory_34 : _GEN_1150; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1152 = 10'h23 == EXMEMALUOut[9:0] ? DMemory_35 : _GEN_1151; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1153 = 10'h24 == EXMEMALUOut[9:0] ? DMemory_36 : _GEN_1152; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1154 = 10'h25 == EXMEMALUOut[9:0] ? DMemory_37 : _GEN_1153; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1155 = 10'h26 == EXMEMALUOut[9:0] ? DMemory_38 : _GEN_1154; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1156 = 10'h27 == EXMEMALUOut[9:0] ? DMemory_39 : _GEN_1155; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1157 = 10'h28 == EXMEMALUOut[9:0] ? DMemory_40 : _GEN_1156; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1158 = 10'h29 == EXMEMALUOut[9:0] ? DMemory_41 : _GEN_1157; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1159 = 10'h2a == EXMEMALUOut[9:0] ? DMemory_42 : _GEN_1158; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1160 = 10'h2b == EXMEMALUOut[9:0] ? DMemory_43 : _GEN_1159; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1161 = 10'h2c == EXMEMALUOut[9:0] ? DMemory_44 : _GEN_1160; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1162 = 10'h2d == EXMEMALUOut[9:0] ? DMemory_45 : _GEN_1161; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1163 = 10'h2e == EXMEMALUOut[9:0] ? DMemory_46 : _GEN_1162; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1164 = 10'h2f == EXMEMALUOut[9:0] ? DMemory_47 : _GEN_1163; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1165 = 10'h30 == EXMEMALUOut[9:0] ? DMemory_48 : _GEN_1164; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1166 = 10'h31 == EXMEMALUOut[9:0] ? DMemory_49 : _GEN_1165; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1167 = 10'h32 == EXMEMALUOut[9:0] ? DMemory_50 : _GEN_1166; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1168 = 10'h33 == EXMEMALUOut[9:0] ? DMemory_51 : _GEN_1167; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1169 = 10'h34 == EXMEMALUOut[9:0] ? DMemory_52 : _GEN_1168; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1170 = 10'h35 == EXMEMALUOut[9:0] ? DMemory_53 : _GEN_1169; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1171 = 10'h36 == EXMEMALUOut[9:0] ? DMemory_54 : _GEN_1170; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1172 = 10'h37 == EXMEMALUOut[9:0] ? DMemory_55 : _GEN_1171; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1173 = 10'h38 == EXMEMALUOut[9:0] ? DMemory_56 : _GEN_1172; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1174 = 10'h39 == EXMEMALUOut[9:0] ? DMemory_57 : _GEN_1173; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1175 = 10'h3a == EXMEMALUOut[9:0] ? DMemory_58 : _GEN_1174; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1176 = 10'h3b == EXMEMALUOut[9:0] ? DMemory_59 : _GEN_1175; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1177 = 10'h3c == EXMEMALUOut[9:0] ? DMemory_60 : _GEN_1176; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1178 = 10'h3d == EXMEMALUOut[9:0] ? DMemory_61 : _GEN_1177; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1179 = 10'h3e == EXMEMALUOut[9:0] ? DMemory_62 : _GEN_1178; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1180 = 10'h3f == EXMEMALUOut[9:0] ? DMemory_63 : _GEN_1179; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1181 = 10'h40 == EXMEMALUOut[9:0] ? DMemory_64 : _GEN_1180; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1182 = 10'h41 == EXMEMALUOut[9:0] ? DMemory_65 : _GEN_1181; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1183 = 10'h42 == EXMEMALUOut[9:0] ? DMemory_66 : _GEN_1182; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1184 = 10'h43 == EXMEMALUOut[9:0] ? DMemory_67 : _GEN_1183; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1185 = 10'h44 == EXMEMALUOut[9:0] ? DMemory_68 : _GEN_1184; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1186 = 10'h45 == EXMEMALUOut[9:0] ? DMemory_69 : _GEN_1185; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1187 = 10'h46 == EXMEMALUOut[9:0] ? DMemory_70 : _GEN_1186; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1188 = 10'h47 == EXMEMALUOut[9:0] ? DMemory_71 : _GEN_1187; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1189 = 10'h48 == EXMEMALUOut[9:0] ? DMemory_72 : _GEN_1188; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1190 = 10'h49 == EXMEMALUOut[9:0] ? DMemory_73 : _GEN_1189; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1191 = 10'h4a == EXMEMALUOut[9:0] ? DMemory_74 : _GEN_1190; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1192 = 10'h4b == EXMEMALUOut[9:0] ? DMemory_75 : _GEN_1191; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1193 = 10'h4c == EXMEMALUOut[9:0] ? DMemory_76 : _GEN_1192; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1194 = 10'h4d == EXMEMALUOut[9:0] ? DMemory_77 : _GEN_1193; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1195 = 10'h4e == EXMEMALUOut[9:0] ? DMemory_78 : _GEN_1194; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1196 = 10'h4f == EXMEMALUOut[9:0] ? DMemory_79 : _GEN_1195; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1197 = 10'h50 == EXMEMALUOut[9:0] ? DMemory_80 : _GEN_1196; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1198 = 10'h51 == EXMEMALUOut[9:0] ? DMemory_81 : _GEN_1197; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1199 = 10'h52 == EXMEMALUOut[9:0] ? DMemory_82 : _GEN_1198; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1200 = 10'h53 == EXMEMALUOut[9:0] ? DMemory_83 : _GEN_1199; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1201 = 10'h54 == EXMEMALUOut[9:0] ? DMemory_84 : _GEN_1200; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1202 = 10'h55 == EXMEMALUOut[9:0] ? DMemory_85 : _GEN_1201; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1203 = 10'h56 == EXMEMALUOut[9:0] ? DMemory_86 : _GEN_1202; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1204 = 10'h57 == EXMEMALUOut[9:0] ? DMemory_87 : _GEN_1203; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1205 = 10'h58 == EXMEMALUOut[9:0] ? DMemory_88 : _GEN_1204; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1206 = 10'h59 == EXMEMALUOut[9:0] ? DMemory_89 : _GEN_1205; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1207 = 10'h5a == EXMEMALUOut[9:0] ? DMemory_90 : _GEN_1206; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1208 = 10'h5b == EXMEMALUOut[9:0] ? DMemory_91 : _GEN_1207; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1209 = 10'h5c == EXMEMALUOut[9:0] ? DMemory_92 : _GEN_1208; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1210 = 10'h5d == EXMEMALUOut[9:0] ? DMemory_93 : _GEN_1209; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1211 = 10'h5e == EXMEMALUOut[9:0] ? DMemory_94 : _GEN_1210; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1212 = 10'h5f == EXMEMALUOut[9:0] ? DMemory_95 : _GEN_1211; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1213 = 10'h60 == EXMEMALUOut[9:0] ? DMemory_96 : _GEN_1212; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1214 = 10'h61 == EXMEMALUOut[9:0] ? DMemory_97 : _GEN_1213; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1215 = 10'h62 == EXMEMALUOut[9:0] ? DMemory_98 : _GEN_1214; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1216 = 10'h63 == EXMEMALUOut[9:0] ? DMemory_99 : _GEN_1215; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1217 = 10'h64 == EXMEMALUOut[9:0] ? DMemory_100 : _GEN_1216; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1218 = 10'h65 == EXMEMALUOut[9:0] ? DMemory_101 : _GEN_1217; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1219 = 10'h66 == EXMEMALUOut[9:0] ? DMemory_102 : _GEN_1218; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1220 = 10'h67 == EXMEMALUOut[9:0] ? DMemory_103 : _GEN_1219; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1221 = 10'h68 == EXMEMALUOut[9:0] ? DMemory_104 : _GEN_1220; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1222 = 10'h69 == EXMEMALUOut[9:0] ? DMemory_105 : _GEN_1221; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1223 = 10'h6a == EXMEMALUOut[9:0] ? DMemory_106 : _GEN_1222; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1224 = 10'h6b == EXMEMALUOut[9:0] ? DMemory_107 : _GEN_1223; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1225 = 10'h6c == EXMEMALUOut[9:0] ? DMemory_108 : _GEN_1224; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1226 = 10'h6d == EXMEMALUOut[9:0] ? DMemory_109 : _GEN_1225; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1227 = 10'h6e == EXMEMALUOut[9:0] ? DMemory_110 : _GEN_1226; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1228 = 10'h6f == EXMEMALUOut[9:0] ? DMemory_111 : _GEN_1227; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1229 = 10'h70 == EXMEMALUOut[9:0] ? DMemory_112 : _GEN_1228; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1230 = 10'h71 == EXMEMALUOut[9:0] ? DMemory_113 : _GEN_1229; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1231 = 10'h72 == EXMEMALUOut[9:0] ? DMemory_114 : _GEN_1230; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1232 = 10'h73 == EXMEMALUOut[9:0] ? DMemory_115 : _GEN_1231; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1233 = 10'h74 == EXMEMALUOut[9:0] ? DMemory_116 : _GEN_1232; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1234 = 10'h75 == EXMEMALUOut[9:0] ? DMemory_117 : _GEN_1233; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1235 = 10'h76 == EXMEMALUOut[9:0] ? DMemory_118 : _GEN_1234; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1236 = 10'h77 == EXMEMALUOut[9:0] ? DMemory_119 : _GEN_1235; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1237 = 10'h78 == EXMEMALUOut[9:0] ? DMemory_120 : _GEN_1236; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1238 = 10'h79 == EXMEMALUOut[9:0] ? DMemory_121 : _GEN_1237; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1239 = 10'h7a == EXMEMALUOut[9:0] ? DMemory_122 : _GEN_1238; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1240 = 10'h7b == EXMEMALUOut[9:0] ? DMemory_123 : _GEN_1239; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1241 = 10'h7c == EXMEMALUOut[9:0] ? DMemory_124 : _GEN_1240; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1242 = 10'h7d == EXMEMALUOut[9:0] ? DMemory_125 : _GEN_1241; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1243 = 10'h7e == EXMEMALUOut[9:0] ? DMemory_126 : _GEN_1242; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1244 = 10'h7f == EXMEMALUOut[9:0] ? DMemory_127 : _GEN_1243; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1245 = 10'h80 == EXMEMALUOut[9:0] ? DMemory_128 : _GEN_1244; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1246 = 10'h81 == EXMEMALUOut[9:0] ? DMemory_129 : _GEN_1245; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1247 = 10'h82 == EXMEMALUOut[9:0] ? DMemory_130 : _GEN_1246; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1248 = 10'h83 == EXMEMALUOut[9:0] ? DMemory_131 : _GEN_1247; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1249 = 10'h84 == EXMEMALUOut[9:0] ? DMemory_132 : _GEN_1248; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1250 = 10'h85 == EXMEMALUOut[9:0] ? DMemory_133 : _GEN_1249; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1251 = 10'h86 == EXMEMALUOut[9:0] ? DMemory_134 : _GEN_1250; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1252 = 10'h87 == EXMEMALUOut[9:0] ? DMemory_135 : _GEN_1251; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1253 = 10'h88 == EXMEMALUOut[9:0] ? DMemory_136 : _GEN_1252; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1254 = 10'h89 == EXMEMALUOut[9:0] ? DMemory_137 : _GEN_1253; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1255 = 10'h8a == EXMEMALUOut[9:0] ? DMemory_138 : _GEN_1254; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1256 = 10'h8b == EXMEMALUOut[9:0] ? DMemory_139 : _GEN_1255; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1257 = 10'h8c == EXMEMALUOut[9:0] ? DMemory_140 : _GEN_1256; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1258 = 10'h8d == EXMEMALUOut[9:0] ? DMemory_141 : _GEN_1257; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1259 = 10'h8e == EXMEMALUOut[9:0] ? DMemory_142 : _GEN_1258; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1260 = 10'h8f == EXMEMALUOut[9:0] ? DMemory_143 : _GEN_1259; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1261 = 10'h90 == EXMEMALUOut[9:0] ? DMemory_144 : _GEN_1260; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1262 = 10'h91 == EXMEMALUOut[9:0] ? DMemory_145 : _GEN_1261; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1263 = 10'h92 == EXMEMALUOut[9:0] ? DMemory_146 : _GEN_1262; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1264 = 10'h93 == EXMEMALUOut[9:0] ? DMemory_147 : _GEN_1263; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1265 = 10'h94 == EXMEMALUOut[9:0] ? DMemory_148 : _GEN_1264; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1266 = 10'h95 == EXMEMALUOut[9:0] ? DMemory_149 : _GEN_1265; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1267 = 10'h96 == EXMEMALUOut[9:0] ? DMemory_150 : _GEN_1266; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1268 = 10'h97 == EXMEMALUOut[9:0] ? DMemory_151 : _GEN_1267; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1269 = 10'h98 == EXMEMALUOut[9:0] ? DMemory_152 : _GEN_1268; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1270 = 10'h99 == EXMEMALUOut[9:0] ? DMemory_153 : _GEN_1269; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1271 = 10'h9a == EXMEMALUOut[9:0] ? DMemory_154 : _GEN_1270; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1272 = 10'h9b == EXMEMALUOut[9:0] ? DMemory_155 : _GEN_1271; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1273 = 10'h9c == EXMEMALUOut[9:0] ? DMemory_156 : _GEN_1272; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1274 = 10'h9d == EXMEMALUOut[9:0] ? DMemory_157 : _GEN_1273; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1275 = 10'h9e == EXMEMALUOut[9:0] ? DMemory_158 : _GEN_1274; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1276 = 10'h9f == EXMEMALUOut[9:0] ? DMemory_159 : _GEN_1275; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1277 = 10'ha0 == EXMEMALUOut[9:0] ? DMemory_160 : _GEN_1276; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1278 = 10'ha1 == EXMEMALUOut[9:0] ? DMemory_161 : _GEN_1277; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1279 = 10'ha2 == EXMEMALUOut[9:0] ? DMemory_162 : _GEN_1278; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1280 = 10'ha3 == EXMEMALUOut[9:0] ? DMemory_163 : _GEN_1279; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1281 = 10'ha4 == EXMEMALUOut[9:0] ? DMemory_164 : _GEN_1280; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1282 = 10'ha5 == EXMEMALUOut[9:0] ? DMemory_165 : _GEN_1281; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1283 = 10'ha6 == EXMEMALUOut[9:0] ? DMemory_166 : _GEN_1282; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1284 = 10'ha7 == EXMEMALUOut[9:0] ? DMemory_167 : _GEN_1283; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1285 = 10'ha8 == EXMEMALUOut[9:0] ? DMemory_168 : _GEN_1284; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1286 = 10'ha9 == EXMEMALUOut[9:0] ? DMemory_169 : _GEN_1285; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1287 = 10'haa == EXMEMALUOut[9:0] ? DMemory_170 : _GEN_1286; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1288 = 10'hab == EXMEMALUOut[9:0] ? DMemory_171 : _GEN_1287; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1289 = 10'hac == EXMEMALUOut[9:0] ? DMemory_172 : _GEN_1288; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1290 = 10'had == EXMEMALUOut[9:0] ? DMemory_173 : _GEN_1289; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1291 = 10'hae == EXMEMALUOut[9:0] ? DMemory_174 : _GEN_1290; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1292 = 10'haf == EXMEMALUOut[9:0] ? DMemory_175 : _GEN_1291; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1293 = 10'hb0 == EXMEMALUOut[9:0] ? DMemory_176 : _GEN_1292; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1294 = 10'hb1 == EXMEMALUOut[9:0] ? DMemory_177 : _GEN_1293; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1295 = 10'hb2 == EXMEMALUOut[9:0] ? DMemory_178 : _GEN_1294; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1296 = 10'hb3 == EXMEMALUOut[9:0] ? DMemory_179 : _GEN_1295; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1297 = 10'hb4 == EXMEMALUOut[9:0] ? DMemory_180 : _GEN_1296; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1298 = 10'hb5 == EXMEMALUOut[9:0] ? DMemory_181 : _GEN_1297; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1299 = 10'hb6 == EXMEMALUOut[9:0] ? DMemory_182 : _GEN_1298; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1300 = 10'hb7 == EXMEMALUOut[9:0] ? DMemory_183 : _GEN_1299; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1301 = 10'hb8 == EXMEMALUOut[9:0] ? DMemory_184 : _GEN_1300; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1302 = 10'hb9 == EXMEMALUOut[9:0] ? DMemory_185 : _GEN_1301; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1303 = 10'hba == EXMEMALUOut[9:0] ? DMemory_186 : _GEN_1302; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1304 = 10'hbb == EXMEMALUOut[9:0] ? DMemory_187 : _GEN_1303; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1305 = 10'hbc == EXMEMALUOut[9:0] ? DMemory_188 : _GEN_1304; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1306 = 10'hbd == EXMEMALUOut[9:0] ? DMemory_189 : _GEN_1305; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1307 = 10'hbe == EXMEMALUOut[9:0] ? DMemory_190 : _GEN_1306; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1308 = 10'hbf == EXMEMALUOut[9:0] ? DMemory_191 : _GEN_1307; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1309 = 10'hc0 == EXMEMALUOut[9:0] ? DMemory_192 : _GEN_1308; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1310 = 10'hc1 == EXMEMALUOut[9:0] ? DMemory_193 : _GEN_1309; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1311 = 10'hc2 == EXMEMALUOut[9:0] ? DMemory_194 : _GEN_1310; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1312 = 10'hc3 == EXMEMALUOut[9:0] ? DMemory_195 : _GEN_1311; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1313 = 10'hc4 == EXMEMALUOut[9:0] ? DMemory_196 : _GEN_1312; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1314 = 10'hc5 == EXMEMALUOut[9:0] ? DMemory_197 : _GEN_1313; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1315 = 10'hc6 == EXMEMALUOut[9:0] ? DMemory_198 : _GEN_1314; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1316 = 10'hc7 == EXMEMALUOut[9:0] ? DMemory_199 : _GEN_1315; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1317 = 10'hc8 == EXMEMALUOut[9:0] ? DMemory_200 : _GEN_1316; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1318 = 10'hc9 == EXMEMALUOut[9:0] ? DMemory_201 : _GEN_1317; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1319 = 10'hca == EXMEMALUOut[9:0] ? DMemory_202 : _GEN_1318; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1320 = 10'hcb == EXMEMALUOut[9:0] ? DMemory_203 : _GEN_1319; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1321 = 10'hcc == EXMEMALUOut[9:0] ? DMemory_204 : _GEN_1320; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1322 = 10'hcd == EXMEMALUOut[9:0] ? DMemory_205 : _GEN_1321; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1323 = 10'hce == EXMEMALUOut[9:0] ? DMemory_206 : _GEN_1322; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1324 = 10'hcf == EXMEMALUOut[9:0] ? DMemory_207 : _GEN_1323; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1325 = 10'hd0 == EXMEMALUOut[9:0] ? DMemory_208 : _GEN_1324; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1326 = 10'hd1 == EXMEMALUOut[9:0] ? DMemory_209 : _GEN_1325; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1327 = 10'hd2 == EXMEMALUOut[9:0] ? DMemory_210 : _GEN_1326; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1328 = 10'hd3 == EXMEMALUOut[9:0] ? DMemory_211 : _GEN_1327; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1329 = 10'hd4 == EXMEMALUOut[9:0] ? DMemory_212 : _GEN_1328; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1330 = 10'hd5 == EXMEMALUOut[9:0] ? DMemory_213 : _GEN_1329; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1331 = 10'hd6 == EXMEMALUOut[9:0] ? DMemory_214 : _GEN_1330; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1332 = 10'hd7 == EXMEMALUOut[9:0] ? DMemory_215 : _GEN_1331; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1333 = 10'hd8 == EXMEMALUOut[9:0] ? DMemory_216 : _GEN_1332; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1334 = 10'hd9 == EXMEMALUOut[9:0] ? DMemory_217 : _GEN_1333; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1335 = 10'hda == EXMEMALUOut[9:0] ? DMemory_218 : _GEN_1334; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1336 = 10'hdb == EXMEMALUOut[9:0] ? DMemory_219 : _GEN_1335; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1337 = 10'hdc == EXMEMALUOut[9:0] ? DMemory_220 : _GEN_1336; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1338 = 10'hdd == EXMEMALUOut[9:0] ? DMemory_221 : _GEN_1337; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1339 = 10'hde == EXMEMALUOut[9:0] ? DMemory_222 : _GEN_1338; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1340 = 10'hdf == EXMEMALUOut[9:0] ? DMemory_223 : _GEN_1339; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1341 = 10'he0 == EXMEMALUOut[9:0] ? DMemory_224 : _GEN_1340; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1342 = 10'he1 == EXMEMALUOut[9:0] ? DMemory_225 : _GEN_1341; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1343 = 10'he2 == EXMEMALUOut[9:0] ? DMemory_226 : _GEN_1342; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1344 = 10'he3 == EXMEMALUOut[9:0] ? DMemory_227 : _GEN_1343; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1345 = 10'he4 == EXMEMALUOut[9:0] ? DMemory_228 : _GEN_1344; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1346 = 10'he5 == EXMEMALUOut[9:0] ? DMemory_229 : _GEN_1345; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1347 = 10'he6 == EXMEMALUOut[9:0] ? DMemory_230 : _GEN_1346; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1348 = 10'he7 == EXMEMALUOut[9:0] ? DMemory_231 : _GEN_1347; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1349 = 10'he8 == EXMEMALUOut[9:0] ? DMemory_232 : _GEN_1348; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1350 = 10'he9 == EXMEMALUOut[9:0] ? DMemory_233 : _GEN_1349; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1351 = 10'hea == EXMEMALUOut[9:0] ? DMemory_234 : _GEN_1350; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1352 = 10'heb == EXMEMALUOut[9:0] ? DMemory_235 : _GEN_1351; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1353 = 10'hec == EXMEMALUOut[9:0] ? DMemory_236 : _GEN_1352; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1354 = 10'hed == EXMEMALUOut[9:0] ? DMemory_237 : _GEN_1353; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1355 = 10'hee == EXMEMALUOut[9:0] ? DMemory_238 : _GEN_1354; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1356 = 10'hef == EXMEMALUOut[9:0] ? DMemory_239 : _GEN_1355; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1357 = 10'hf0 == EXMEMALUOut[9:0] ? DMemory_240 : _GEN_1356; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1358 = 10'hf1 == EXMEMALUOut[9:0] ? DMemory_241 : _GEN_1357; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1359 = 10'hf2 == EXMEMALUOut[9:0] ? DMemory_242 : _GEN_1358; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1360 = 10'hf3 == EXMEMALUOut[9:0] ? DMemory_243 : _GEN_1359; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1361 = 10'hf4 == EXMEMALUOut[9:0] ? DMemory_244 : _GEN_1360; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1362 = 10'hf5 == EXMEMALUOut[9:0] ? DMemory_245 : _GEN_1361; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1363 = 10'hf6 == EXMEMALUOut[9:0] ? DMemory_246 : _GEN_1362; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1364 = 10'hf7 == EXMEMALUOut[9:0] ? DMemory_247 : _GEN_1363; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1365 = 10'hf8 == EXMEMALUOut[9:0] ? DMemory_248 : _GEN_1364; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1366 = 10'hf9 == EXMEMALUOut[9:0] ? DMemory_249 : _GEN_1365; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1367 = 10'hfa == EXMEMALUOut[9:0] ? DMemory_250 : _GEN_1366; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1368 = 10'hfb == EXMEMALUOut[9:0] ? DMemory_251 : _GEN_1367; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1369 = 10'hfc == EXMEMALUOut[9:0] ? DMemory_252 : _GEN_1368; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1370 = 10'hfd == EXMEMALUOut[9:0] ? DMemory_253 : _GEN_1369; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1371 = 10'hfe == EXMEMALUOut[9:0] ? DMemory_254 : _GEN_1370; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1372 = 10'hff == EXMEMALUOut[9:0] ? DMemory_255 : _GEN_1371; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1373 = 10'h100 == EXMEMALUOut[9:0] ? DMemory_256 : _GEN_1372; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1374 = 10'h101 == EXMEMALUOut[9:0] ? DMemory_257 : _GEN_1373; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1375 = 10'h102 == EXMEMALUOut[9:0] ? DMemory_258 : _GEN_1374; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1376 = 10'h103 == EXMEMALUOut[9:0] ? DMemory_259 : _GEN_1375; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1377 = 10'h104 == EXMEMALUOut[9:0] ? DMemory_260 : _GEN_1376; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1378 = 10'h105 == EXMEMALUOut[9:0] ? DMemory_261 : _GEN_1377; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1379 = 10'h106 == EXMEMALUOut[9:0] ? DMemory_262 : _GEN_1378; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1380 = 10'h107 == EXMEMALUOut[9:0] ? DMemory_263 : _GEN_1379; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1381 = 10'h108 == EXMEMALUOut[9:0] ? DMemory_264 : _GEN_1380; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1382 = 10'h109 == EXMEMALUOut[9:0] ? DMemory_265 : _GEN_1381; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1383 = 10'h10a == EXMEMALUOut[9:0] ? DMemory_266 : _GEN_1382; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1384 = 10'h10b == EXMEMALUOut[9:0] ? DMemory_267 : _GEN_1383; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1385 = 10'h10c == EXMEMALUOut[9:0] ? DMemory_268 : _GEN_1384; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1386 = 10'h10d == EXMEMALUOut[9:0] ? DMemory_269 : _GEN_1385; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1387 = 10'h10e == EXMEMALUOut[9:0] ? DMemory_270 : _GEN_1386; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1388 = 10'h10f == EXMEMALUOut[9:0] ? DMemory_271 : _GEN_1387; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1389 = 10'h110 == EXMEMALUOut[9:0] ? DMemory_272 : _GEN_1388; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1390 = 10'h111 == EXMEMALUOut[9:0] ? DMemory_273 : _GEN_1389; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1391 = 10'h112 == EXMEMALUOut[9:0] ? DMemory_274 : _GEN_1390; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1392 = 10'h113 == EXMEMALUOut[9:0] ? DMemory_275 : _GEN_1391; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1393 = 10'h114 == EXMEMALUOut[9:0] ? DMemory_276 : _GEN_1392; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1394 = 10'h115 == EXMEMALUOut[9:0] ? DMemory_277 : _GEN_1393; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1395 = 10'h116 == EXMEMALUOut[9:0] ? DMemory_278 : _GEN_1394; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1396 = 10'h117 == EXMEMALUOut[9:0] ? DMemory_279 : _GEN_1395; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1397 = 10'h118 == EXMEMALUOut[9:0] ? DMemory_280 : _GEN_1396; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1398 = 10'h119 == EXMEMALUOut[9:0] ? DMemory_281 : _GEN_1397; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1399 = 10'h11a == EXMEMALUOut[9:0] ? DMemory_282 : _GEN_1398; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1400 = 10'h11b == EXMEMALUOut[9:0] ? DMemory_283 : _GEN_1399; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1401 = 10'h11c == EXMEMALUOut[9:0] ? DMemory_284 : _GEN_1400; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1402 = 10'h11d == EXMEMALUOut[9:0] ? DMemory_285 : _GEN_1401; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1403 = 10'h11e == EXMEMALUOut[9:0] ? DMemory_286 : _GEN_1402; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1404 = 10'h11f == EXMEMALUOut[9:0] ? DMemory_287 : _GEN_1403; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1405 = 10'h120 == EXMEMALUOut[9:0] ? DMemory_288 : _GEN_1404; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1406 = 10'h121 == EXMEMALUOut[9:0] ? DMemory_289 : _GEN_1405; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1407 = 10'h122 == EXMEMALUOut[9:0] ? DMemory_290 : _GEN_1406; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1408 = 10'h123 == EXMEMALUOut[9:0] ? DMemory_291 : _GEN_1407; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1409 = 10'h124 == EXMEMALUOut[9:0] ? DMemory_292 : _GEN_1408; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1410 = 10'h125 == EXMEMALUOut[9:0] ? DMemory_293 : _GEN_1409; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1411 = 10'h126 == EXMEMALUOut[9:0] ? DMemory_294 : _GEN_1410; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1412 = 10'h127 == EXMEMALUOut[9:0] ? DMemory_295 : _GEN_1411; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1413 = 10'h128 == EXMEMALUOut[9:0] ? DMemory_296 : _GEN_1412; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1414 = 10'h129 == EXMEMALUOut[9:0] ? DMemory_297 : _GEN_1413; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1415 = 10'h12a == EXMEMALUOut[9:0] ? DMemory_298 : _GEN_1414; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1416 = 10'h12b == EXMEMALUOut[9:0] ? DMemory_299 : _GEN_1415; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1417 = 10'h12c == EXMEMALUOut[9:0] ? DMemory_300 : _GEN_1416; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1418 = 10'h12d == EXMEMALUOut[9:0] ? DMemory_301 : _GEN_1417; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1419 = 10'h12e == EXMEMALUOut[9:0] ? DMemory_302 : _GEN_1418; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1420 = 10'h12f == EXMEMALUOut[9:0] ? DMemory_303 : _GEN_1419; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1421 = 10'h130 == EXMEMALUOut[9:0] ? DMemory_304 : _GEN_1420; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1422 = 10'h131 == EXMEMALUOut[9:0] ? DMemory_305 : _GEN_1421; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1423 = 10'h132 == EXMEMALUOut[9:0] ? DMemory_306 : _GEN_1422; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1424 = 10'h133 == EXMEMALUOut[9:0] ? DMemory_307 : _GEN_1423; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1425 = 10'h134 == EXMEMALUOut[9:0] ? DMemory_308 : _GEN_1424; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1426 = 10'h135 == EXMEMALUOut[9:0] ? DMemory_309 : _GEN_1425; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1427 = 10'h136 == EXMEMALUOut[9:0] ? DMemory_310 : _GEN_1426; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1428 = 10'h137 == EXMEMALUOut[9:0] ? DMemory_311 : _GEN_1427; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1429 = 10'h138 == EXMEMALUOut[9:0] ? DMemory_312 : _GEN_1428; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1430 = 10'h139 == EXMEMALUOut[9:0] ? DMemory_313 : _GEN_1429; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1431 = 10'h13a == EXMEMALUOut[9:0] ? DMemory_314 : _GEN_1430; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1432 = 10'h13b == EXMEMALUOut[9:0] ? DMemory_315 : _GEN_1431; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1433 = 10'h13c == EXMEMALUOut[9:0] ? DMemory_316 : _GEN_1432; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1434 = 10'h13d == EXMEMALUOut[9:0] ? DMemory_317 : _GEN_1433; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1435 = 10'h13e == EXMEMALUOut[9:0] ? DMemory_318 : _GEN_1434; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1436 = 10'h13f == EXMEMALUOut[9:0] ? DMemory_319 : _GEN_1435; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1437 = 10'h140 == EXMEMALUOut[9:0] ? DMemory_320 : _GEN_1436; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1438 = 10'h141 == EXMEMALUOut[9:0] ? DMemory_321 : _GEN_1437; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1439 = 10'h142 == EXMEMALUOut[9:0] ? DMemory_322 : _GEN_1438; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1440 = 10'h143 == EXMEMALUOut[9:0] ? DMemory_323 : _GEN_1439; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1441 = 10'h144 == EXMEMALUOut[9:0] ? DMemory_324 : _GEN_1440; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1442 = 10'h145 == EXMEMALUOut[9:0] ? DMemory_325 : _GEN_1441; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1443 = 10'h146 == EXMEMALUOut[9:0] ? DMemory_326 : _GEN_1442; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1444 = 10'h147 == EXMEMALUOut[9:0] ? DMemory_327 : _GEN_1443; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1445 = 10'h148 == EXMEMALUOut[9:0] ? DMemory_328 : _GEN_1444; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1446 = 10'h149 == EXMEMALUOut[9:0] ? DMemory_329 : _GEN_1445; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1447 = 10'h14a == EXMEMALUOut[9:0] ? DMemory_330 : _GEN_1446; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1448 = 10'h14b == EXMEMALUOut[9:0] ? DMemory_331 : _GEN_1447; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1449 = 10'h14c == EXMEMALUOut[9:0] ? DMemory_332 : _GEN_1448; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1450 = 10'h14d == EXMEMALUOut[9:0] ? DMemory_333 : _GEN_1449; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1451 = 10'h14e == EXMEMALUOut[9:0] ? DMemory_334 : _GEN_1450; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1452 = 10'h14f == EXMEMALUOut[9:0] ? DMemory_335 : _GEN_1451; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1453 = 10'h150 == EXMEMALUOut[9:0] ? DMemory_336 : _GEN_1452; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1454 = 10'h151 == EXMEMALUOut[9:0] ? DMemory_337 : _GEN_1453; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1455 = 10'h152 == EXMEMALUOut[9:0] ? DMemory_338 : _GEN_1454; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1456 = 10'h153 == EXMEMALUOut[9:0] ? DMemory_339 : _GEN_1455; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1457 = 10'h154 == EXMEMALUOut[9:0] ? DMemory_340 : _GEN_1456; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1458 = 10'h155 == EXMEMALUOut[9:0] ? DMemory_341 : _GEN_1457; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1459 = 10'h156 == EXMEMALUOut[9:0] ? DMemory_342 : _GEN_1458; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1460 = 10'h157 == EXMEMALUOut[9:0] ? DMemory_343 : _GEN_1459; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1461 = 10'h158 == EXMEMALUOut[9:0] ? DMemory_344 : _GEN_1460; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1462 = 10'h159 == EXMEMALUOut[9:0] ? DMemory_345 : _GEN_1461; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1463 = 10'h15a == EXMEMALUOut[9:0] ? DMemory_346 : _GEN_1462; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1464 = 10'h15b == EXMEMALUOut[9:0] ? DMemory_347 : _GEN_1463; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1465 = 10'h15c == EXMEMALUOut[9:0] ? DMemory_348 : _GEN_1464; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1466 = 10'h15d == EXMEMALUOut[9:0] ? DMemory_349 : _GEN_1465; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1467 = 10'h15e == EXMEMALUOut[9:0] ? DMemory_350 : _GEN_1466; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1468 = 10'h15f == EXMEMALUOut[9:0] ? DMemory_351 : _GEN_1467; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1469 = 10'h160 == EXMEMALUOut[9:0] ? DMemory_352 : _GEN_1468; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1470 = 10'h161 == EXMEMALUOut[9:0] ? DMemory_353 : _GEN_1469; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1471 = 10'h162 == EXMEMALUOut[9:0] ? DMemory_354 : _GEN_1470; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1472 = 10'h163 == EXMEMALUOut[9:0] ? DMemory_355 : _GEN_1471; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1473 = 10'h164 == EXMEMALUOut[9:0] ? DMemory_356 : _GEN_1472; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1474 = 10'h165 == EXMEMALUOut[9:0] ? DMemory_357 : _GEN_1473; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1475 = 10'h166 == EXMEMALUOut[9:0] ? DMemory_358 : _GEN_1474; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1476 = 10'h167 == EXMEMALUOut[9:0] ? DMemory_359 : _GEN_1475; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1477 = 10'h168 == EXMEMALUOut[9:0] ? DMemory_360 : _GEN_1476; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1478 = 10'h169 == EXMEMALUOut[9:0] ? DMemory_361 : _GEN_1477; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1479 = 10'h16a == EXMEMALUOut[9:0] ? DMemory_362 : _GEN_1478; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1480 = 10'h16b == EXMEMALUOut[9:0] ? DMemory_363 : _GEN_1479; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1481 = 10'h16c == EXMEMALUOut[9:0] ? DMemory_364 : _GEN_1480; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1482 = 10'h16d == EXMEMALUOut[9:0] ? DMemory_365 : _GEN_1481; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1483 = 10'h16e == EXMEMALUOut[9:0] ? DMemory_366 : _GEN_1482; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1484 = 10'h16f == EXMEMALUOut[9:0] ? DMemory_367 : _GEN_1483; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1485 = 10'h170 == EXMEMALUOut[9:0] ? DMemory_368 : _GEN_1484; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1486 = 10'h171 == EXMEMALUOut[9:0] ? DMemory_369 : _GEN_1485; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1487 = 10'h172 == EXMEMALUOut[9:0] ? DMemory_370 : _GEN_1486; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1488 = 10'h173 == EXMEMALUOut[9:0] ? DMemory_371 : _GEN_1487; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1489 = 10'h174 == EXMEMALUOut[9:0] ? DMemory_372 : _GEN_1488; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1490 = 10'h175 == EXMEMALUOut[9:0] ? DMemory_373 : _GEN_1489; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1491 = 10'h176 == EXMEMALUOut[9:0] ? DMemory_374 : _GEN_1490; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1492 = 10'h177 == EXMEMALUOut[9:0] ? DMemory_375 : _GEN_1491; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1493 = 10'h178 == EXMEMALUOut[9:0] ? DMemory_376 : _GEN_1492; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1494 = 10'h179 == EXMEMALUOut[9:0] ? DMemory_377 : _GEN_1493; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1495 = 10'h17a == EXMEMALUOut[9:0] ? DMemory_378 : _GEN_1494; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1496 = 10'h17b == EXMEMALUOut[9:0] ? DMemory_379 : _GEN_1495; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1497 = 10'h17c == EXMEMALUOut[9:0] ? DMemory_380 : _GEN_1496; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1498 = 10'h17d == EXMEMALUOut[9:0] ? DMemory_381 : _GEN_1497; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1499 = 10'h17e == EXMEMALUOut[9:0] ? DMemory_382 : _GEN_1498; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1500 = 10'h17f == EXMEMALUOut[9:0] ? DMemory_383 : _GEN_1499; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1501 = 10'h180 == EXMEMALUOut[9:0] ? DMemory_384 : _GEN_1500; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1502 = 10'h181 == EXMEMALUOut[9:0] ? DMemory_385 : _GEN_1501; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1503 = 10'h182 == EXMEMALUOut[9:0] ? DMemory_386 : _GEN_1502; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1504 = 10'h183 == EXMEMALUOut[9:0] ? DMemory_387 : _GEN_1503; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1505 = 10'h184 == EXMEMALUOut[9:0] ? DMemory_388 : _GEN_1504; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1506 = 10'h185 == EXMEMALUOut[9:0] ? DMemory_389 : _GEN_1505; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1507 = 10'h186 == EXMEMALUOut[9:0] ? DMemory_390 : _GEN_1506; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1508 = 10'h187 == EXMEMALUOut[9:0] ? DMemory_391 : _GEN_1507; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1509 = 10'h188 == EXMEMALUOut[9:0] ? DMemory_392 : _GEN_1508; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1510 = 10'h189 == EXMEMALUOut[9:0] ? DMemory_393 : _GEN_1509; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1511 = 10'h18a == EXMEMALUOut[9:0] ? DMemory_394 : _GEN_1510; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1512 = 10'h18b == EXMEMALUOut[9:0] ? DMemory_395 : _GEN_1511; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1513 = 10'h18c == EXMEMALUOut[9:0] ? DMemory_396 : _GEN_1512; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1514 = 10'h18d == EXMEMALUOut[9:0] ? DMemory_397 : _GEN_1513; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1515 = 10'h18e == EXMEMALUOut[9:0] ? DMemory_398 : _GEN_1514; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1516 = 10'h18f == EXMEMALUOut[9:0] ? DMemory_399 : _GEN_1515; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1517 = 10'h190 == EXMEMALUOut[9:0] ? DMemory_400 : _GEN_1516; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1518 = 10'h191 == EXMEMALUOut[9:0] ? DMemory_401 : _GEN_1517; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1519 = 10'h192 == EXMEMALUOut[9:0] ? DMemory_402 : _GEN_1518; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1520 = 10'h193 == EXMEMALUOut[9:0] ? DMemory_403 : _GEN_1519; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1521 = 10'h194 == EXMEMALUOut[9:0] ? DMemory_404 : _GEN_1520; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1522 = 10'h195 == EXMEMALUOut[9:0] ? DMemory_405 : _GEN_1521; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1523 = 10'h196 == EXMEMALUOut[9:0] ? DMemory_406 : _GEN_1522; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1524 = 10'h197 == EXMEMALUOut[9:0] ? DMemory_407 : _GEN_1523; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1525 = 10'h198 == EXMEMALUOut[9:0] ? DMemory_408 : _GEN_1524; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1526 = 10'h199 == EXMEMALUOut[9:0] ? DMemory_409 : _GEN_1525; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1527 = 10'h19a == EXMEMALUOut[9:0] ? DMemory_410 : _GEN_1526; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1528 = 10'h19b == EXMEMALUOut[9:0] ? DMemory_411 : _GEN_1527; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1529 = 10'h19c == EXMEMALUOut[9:0] ? DMemory_412 : _GEN_1528; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1530 = 10'h19d == EXMEMALUOut[9:0] ? DMemory_413 : _GEN_1529; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1531 = 10'h19e == EXMEMALUOut[9:0] ? DMemory_414 : _GEN_1530; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1532 = 10'h19f == EXMEMALUOut[9:0] ? DMemory_415 : _GEN_1531; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1533 = 10'h1a0 == EXMEMALUOut[9:0] ? DMemory_416 : _GEN_1532; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1534 = 10'h1a1 == EXMEMALUOut[9:0] ? DMemory_417 : _GEN_1533; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1535 = 10'h1a2 == EXMEMALUOut[9:0] ? DMemory_418 : _GEN_1534; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1536 = 10'h1a3 == EXMEMALUOut[9:0] ? DMemory_419 : _GEN_1535; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1537 = 10'h1a4 == EXMEMALUOut[9:0] ? DMemory_420 : _GEN_1536; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1538 = 10'h1a5 == EXMEMALUOut[9:0] ? DMemory_421 : _GEN_1537; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1539 = 10'h1a6 == EXMEMALUOut[9:0] ? DMemory_422 : _GEN_1538; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1540 = 10'h1a7 == EXMEMALUOut[9:0] ? DMemory_423 : _GEN_1539; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1541 = 10'h1a8 == EXMEMALUOut[9:0] ? DMemory_424 : _GEN_1540; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1542 = 10'h1a9 == EXMEMALUOut[9:0] ? DMemory_425 : _GEN_1541; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1543 = 10'h1aa == EXMEMALUOut[9:0] ? DMemory_426 : _GEN_1542; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1544 = 10'h1ab == EXMEMALUOut[9:0] ? DMemory_427 : _GEN_1543; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1545 = 10'h1ac == EXMEMALUOut[9:0] ? DMemory_428 : _GEN_1544; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1546 = 10'h1ad == EXMEMALUOut[9:0] ? DMemory_429 : _GEN_1545; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1547 = 10'h1ae == EXMEMALUOut[9:0] ? DMemory_430 : _GEN_1546; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1548 = 10'h1af == EXMEMALUOut[9:0] ? DMemory_431 : _GEN_1547; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1549 = 10'h1b0 == EXMEMALUOut[9:0] ? DMemory_432 : _GEN_1548; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1550 = 10'h1b1 == EXMEMALUOut[9:0] ? DMemory_433 : _GEN_1549; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1551 = 10'h1b2 == EXMEMALUOut[9:0] ? DMemory_434 : _GEN_1550; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1552 = 10'h1b3 == EXMEMALUOut[9:0] ? DMemory_435 : _GEN_1551; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1553 = 10'h1b4 == EXMEMALUOut[9:0] ? DMemory_436 : _GEN_1552; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1554 = 10'h1b5 == EXMEMALUOut[9:0] ? DMemory_437 : _GEN_1553; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1555 = 10'h1b6 == EXMEMALUOut[9:0] ? DMemory_438 : _GEN_1554; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1556 = 10'h1b7 == EXMEMALUOut[9:0] ? DMemory_439 : _GEN_1555; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1557 = 10'h1b8 == EXMEMALUOut[9:0] ? DMemory_440 : _GEN_1556; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1558 = 10'h1b9 == EXMEMALUOut[9:0] ? DMemory_441 : _GEN_1557; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1559 = 10'h1ba == EXMEMALUOut[9:0] ? DMemory_442 : _GEN_1558; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1560 = 10'h1bb == EXMEMALUOut[9:0] ? DMemory_443 : _GEN_1559; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1561 = 10'h1bc == EXMEMALUOut[9:0] ? DMemory_444 : _GEN_1560; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1562 = 10'h1bd == EXMEMALUOut[9:0] ? DMemory_445 : _GEN_1561; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1563 = 10'h1be == EXMEMALUOut[9:0] ? DMemory_446 : _GEN_1562; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1564 = 10'h1bf == EXMEMALUOut[9:0] ? DMemory_447 : _GEN_1563; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1565 = 10'h1c0 == EXMEMALUOut[9:0] ? DMemory_448 : _GEN_1564; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1566 = 10'h1c1 == EXMEMALUOut[9:0] ? DMemory_449 : _GEN_1565; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1567 = 10'h1c2 == EXMEMALUOut[9:0] ? DMemory_450 : _GEN_1566; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1568 = 10'h1c3 == EXMEMALUOut[9:0] ? DMemory_451 : _GEN_1567; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1569 = 10'h1c4 == EXMEMALUOut[9:0] ? DMemory_452 : _GEN_1568; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1570 = 10'h1c5 == EXMEMALUOut[9:0] ? DMemory_453 : _GEN_1569; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1571 = 10'h1c6 == EXMEMALUOut[9:0] ? DMemory_454 : _GEN_1570; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1572 = 10'h1c7 == EXMEMALUOut[9:0] ? DMemory_455 : _GEN_1571; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1573 = 10'h1c8 == EXMEMALUOut[9:0] ? DMemory_456 : _GEN_1572; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1574 = 10'h1c9 == EXMEMALUOut[9:0] ? DMemory_457 : _GEN_1573; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1575 = 10'h1ca == EXMEMALUOut[9:0] ? DMemory_458 : _GEN_1574; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1576 = 10'h1cb == EXMEMALUOut[9:0] ? DMemory_459 : _GEN_1575; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1577 = 10'h1cc == EXMEMALUOut[9:0] ? DMemory_460 : _GEN_1576; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1578 = 10'h1cd == EXMEMALUOut[9:0] ? DMemory_461 : _GEN_1577; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1579 = 10'h1ce == EXMEMALUOut[9:0] ? DMemory_462 : _GEN_1578; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1580 = 10'h1cf == EXMEMALUOut[9:0] ? DMemory_463 : _GEN_1579; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1581 = 10'h1d0 == EXMEMALUOut[9:0] ? DMemory_464 : _GEN_1580; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1582 = 10'h1d1 == EXMEMALUOut[9:0] ? DMemory_465 : _GEN_1581; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1583 = 10'h1d2 == EXMEMALUOut[9:0] ? DMemory_466 : _GEN_1582; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1584 = 10'h1d3 == EXMEMALUOut[9:0] ? DMemory_467 : _GEN_1583; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1585 = 10'h1d4 == EXMEMALUOut[9:0] ? DMemory_468 : _GEN_1584; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1586 = 10'h1d5 == EXMEMALUOut[9:0] ? DMemory_469 : _GEN_1585; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1587 = 10'h1d6 == EXMEMALUOut[9:0] ? DMemory_470 : _GEN_1586; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1588 = 10'h1d7 == EXMEMALUOut[9:0] ? DMemory_471 : _GEN_1587; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1589 = 10'h1d8 == EXMEMALUOut[9:0] ? DMemory_472 : _GEN_1588; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1590 = 10'h1d9 == EXMEMALUOut[9:0] ? DMemory_473 : _GEN_1589; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1591 = 10'h1da == EXMEMALUOut[9:0] ? DMemory_474 : _GEN_1590; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1592 = 10'h1db == EXMEMALUOut[9:0] ? DMemory_475 : _GEN_1591; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1593 = 10'h1dc == EXMEMALUOut[9:0] ? DMemory_476 : _GEN_1592; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1594 = 10'h1dd == EXMEMALUOut[9:0] ? DMemory_477 : _GEN_1593; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1595 = 10'h1de == EXMEMALUOut[9:0] ? DMemory_478 : _GEN_1594; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1596 = 10'h1df == EXMEMALUOut[9:0] ? DMemory_479 : _GEN_1595; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1597 = 10'h1e0 == EXMEMALUOut[9:0] ? DMemory_480 : _GEN_1596; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1598 = 10'h1e1 == EXMEMALUOut[9:0] ? DMemory_481 : _GEN_1597; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1599 = 10'h1e2 == EXMEMALUOut[9:0] ? DMemory_482 : _GEN_1598; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1600 = 10'h1e3 == EXMEMALUOut[9:0] ? DMemory_483 : _GEN_1599; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1601 = 10'h1e4 == EXMEMALUOut[9:0] ? DMemory_484 : _GEN_1600; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1602 = 10'h1e5 == EXMEMALUOut[9:0] ? DMemory_485 : _GEN_1601; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1603 = 10'h1e6 == EXMEMALUOut[9:0] ? DMemory_486 : _GEN_1602; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1604 = 10'h1e7 == EXMEMALUOut[9:0] ? DMemory_487 : _GEN_1603; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1605 = 10'h1e8 == EXMEMALUOut[9:0] ? DMemory_488 : _GEN_1604; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1606 = 10'h1e9 == EXMEMALUOut[9:0] ? DMemory_489 : _GEN_1605; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1607 = 10'h1ea == EXMEMALUOut[9:0] ? DMemory_490 : _GEN_1606; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1608 = 10'h1eb == EXMEMALUOut[9:0] ? DMemory_491 : _GEN_1607; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1609 = 10'h1ec == EXMEMALUOut[9:0] ? DMemory_492 : _GEN_1608; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1610 = 10'h1ed == EXMEMALUOut[9:0] ? DMemory_493 : _GEN_1609; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1611 = 10'h1ee == EXMEMALUOut[9:0] ? DMemory_494 : _GEN_1610; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1612 = 10'h1ef == EXMEMALUOut[9:0] ? DMemory_495 : _GEN_1611; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1613 = 10'h1f0 == EXMEMALUOut[9:0] ? DMemory_496 : _GEN_1612; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1614 = 10'h1f1 == EXMEMALUOut[9:0] ? DMemory_497 : _GEN_1613; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1615 = 10'h1f2 == EXMEMALUOut[9:0] ? DMemory_498 : _GEN_1614; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1616 = 10'h1f3 == EXMEMALUOut[9:0] ? DMemory_499 : _GEN_1615; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1617 = 10'h1f4 == EXMEMALUOut[9:0] ? DMemory_500 : _GEN_1616; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1618 = 10'h1f5 == EXMEMALUOut[9:0] ? DMemory_501 : _GEN_1617; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1619 = 10'h1f6 == EXMEMALUOut[9:0] ? DMemory_502 : _GEN_1618; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1620 = 10'h1f7 == EXMEMALUOut[9:0] ? DMemory_503 : _GEN_1619; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1621 = 10'h1f8 == EXMEMALUOut[9:0] ? DMemory_504 : _GEN_1620; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1622 = 10'h1f9 == EXMEMALUOut[9:0] ? DMemory_505 : _GEN_1621; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1623 = 10'h1fa == EXMEMALUOut[9:0] ? DMemory_506 : _GEN_1622; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1624 = 10'h1fb == EXMEMALUOut[9:0] ? DMemory_507 : _GEN_1623; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1625 = 10'h1fc == EXMEMALUOut[9:0] ? DMemory_508 : _GEN_1624; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1626 = 10'h1fd == EXMEMALUOut[9:0] ? DMemory_509 : _GEN_1625; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1627 = 10'h1fe == EXMEMALUOut[9:0] ? DMemory_510 : _GEN_1626; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1628 = 10'h1ff == EXMEMALUOut[9:0] ? DMemory_511 : _GEN_1627; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1629 = 10'h200 == EXMEMALUOut[9:0] ? DMemory_512 : _GEN_1628; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1630 = 10'h201 == EXMEMALUOut[9:0] ? DMemory_513 : _GEN_1629; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1631 = 10'h202 == EXMEMALUOut[9:0] ? DMemory_514 : _GEN_1630; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1632 = 10'h203 == EXMEMALUOut[9:0] ? DMemory_515 : _GEN_1631; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1633 = 10'h204 == EXMEMALUOut[9:0] ? DMemory_516 : _GEN_1632; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1634 = 10'h205 == EXMEMALUOut[9:0] ? DMemory_517 : _GEN_1633; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1635 = 10'h206 == EXMEMALUOut[9:0] ? DMemory_518 : _GEN_1634; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1636 = 10'h207 == EXMEMALUOut[9:0] ? DMemory_519 : _GEN_1635; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1637 = 10'h208 == EXMEMALUOut[9:0] ? DMemory_520 : _GEN_1636; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1638 = 10'h209 == EXMEMALUOut[9:0] ? DMemory_521 : _GEN_1637; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1639 = 10'h20a == EXMEMALUOut[9:0] ? DMemory_522 : _GEN_1638; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1640 = 10'h20b == EXMEMALUOut[9:0] ? DMemory_523 : _GEN_1639; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1641 = 10'h20c == EXMEMALUOut[9:0] ? DMemory_524 : _GEN_1640; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1642 = 10'h20d == EXMEMALUOut[9:0] ? DMemory_525 : _GEN_1641; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1643 = 10'h20e == EXMEMALUOut[9:0] ? DMemory_526 : _GEN_1642; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1644 = 10'h20f == EXMEMALUOut[9:0] ? DMemory_527 : _GEN_1643; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1645 = 10'h210 == EXMEMALUOut[9:0] ? DMemory_528 : _GEN_1644; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1646 = 10'h211 == EXMEMALUOut[9:0] ? DMemory_529 : _GEN_1645; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1647 = 10'h212 == EXMEMALUOut[9:0] ? DMemory_530 : _GEN_1646; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1648 = 10'h213 == EXMEMALUOut[9:0] ? DMemory_531 : _GEN_1647; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1649 = 10'h214 == EXMEMALUOut[9:0] ? DMemory_532 : _GEN_1648; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1650 = 10'h215 == EXMEMALUOut[9:0] ? DMemory_533 : _GEN_1649; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1651 = 10'h216 == EXMEMALUOut[9:0] ? DMemory_534 : _GEN_1650; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1652 = 10'h217 == EXMEMALUOut[9:0] ? DMemory_535 : _GEN_1651; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1653 = 10'h218 == EXMEMALUOut[9:0] ? DMemory_536 : _GEN_1652; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1654 = 10'h219 == EXMEMALUOut[9:0] ? DMemory_537 : _GEN_1653; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1655 = 10'h21a == EXMEMALUOut[9:0] ? DMemory_538 : _GEN_1654; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1656 = 10'h21b == EXMEMALUOut[9:0] ? DMemory_539 : _GEN_1655; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1657 = 10'h21c == EXMEMALUOut[9:0] ? DMemory_540 : _GEN_1656; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1658 = 10'h21d == EXMEMALUOut[9:0] ? DMemory_541 : _GEN_1657; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1659 = 10'h21e == EXMEMALUOut[9:0] ? DMemory_542 : _GEN_1658; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1660 = 10'h21f == EXMEMALUOut[9:0] ? DMemory_543 : _GEN_1659; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1661 = 10'h220 == EXMEMALUOut[9:0] ? DMemory_544 : _GEN_1660; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1662 = 10'h221 == EXMEMALUOut[9:0] ? DMemory_545 : _GEN_1661; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1663 = 10'h222 == EXMEMALUOut[9:0] ? DMemory_546 : _GEN_1662; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1664 = 10'h223 == EXMEMALUOut[9:0] ? DMemory_547 : _GEN_1663; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1665 = 10'h224 == EXMEMALUOut[9:0] ? DMemory_548 : _GEN_1664; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1666 = 10'h225 == EXMEMALUOut[9:0] ? DMemory_549 : _GEN_1665; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1667 = 10'h226 == EXMEMALUOut[9:0] ? DMemory_550 : _GEN_1666; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1668 = 10'h227 == EXMEMALUOut[9:0] ? DMemory_551 : _GEN_1667; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1669 = 10'h228 == EXMEMALUOut[9:0] ? DMemory_552 : _GEN_1668; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1670 = 10'h229 == EXMEMALUOut[9:0] ? DMemory_553 : _GEN_1669; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1671 = 10'h22a == EXMEMALUOut[9:0] ? DMemory_554 : _GEN_1670; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1672 = 10'h22b == EXMEMALUOut[9:0] ? DMemory_555 : _GEN_1671; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1673 = 10'h22c == EXMEMALUOut[9:0] ? DMemory_556 : _GEN_1672; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1674 = 10'h22d == EXMEMALUOut[9:0] ? DMemory_557 : _GEN_1673; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1675 = 10'h22e == EXMEMALUOut[9:0] ? DMemory_558 : _GEN_1674; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1676 = 10'h22f == EXMEMALUOut[9:0] ? DMemory_559 : _GEN_1675; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1677 = 10'h230 == EXMEMALUOut[9:0] ? DMemory_560 : _GEN_1676; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1678 = 10'h231 == EXMEMALUOut[9:0] ? DMemory_561 : _GEN_1677; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1679 = 10'h232 == EXMEMALUOut[9:0] ? DMemory_562 : _GEN_1678; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1680 = 10'h233 == EXMEMALUOut[9:0] ? DMemory_563 : _GEN_1679; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1681 = 10'h234 == EXMEMALUOut[9:0] ? DMemory_564 : _GEN_1680; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1682 = 10'h235 == EXMEMALUOut[9:0] ? DMemory_565 : _GEN_1681; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1683 = 10'h236 == EXMEMALUOut[9:0] ? DMemory_566 : _GEN_1682; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1684 = 10'h237 == EXMEMALUOut[9:0] ? DMemory_567 : _GEN_1683; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1685 = 10'h238 == EXMEMALUOut[9:0] ? DMemory_568 : _GEN_1684; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1686 = 10'h239 == EXMEMALUOut[9:0] ? DMemory_569 : _GEN_1685; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1687 = 10'h23a == EXMEMALUOut[9:0] ? DMemory_570 : _GEN_1686; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1688 = 10'h23b == EXMEMALUOut[9:0] ? DMemory_571 : _GEN_1687; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1689 = 10'h23c == EXMEMALUOut[9:0] ? DMemory_572 : _GEN_1688; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1690 = 10'h23d == EXMEMALUOut[9:0] ? DMemory_573 : _GEN_1689; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1691 = 10'h23e == EXMEMALUOut[9:0] ? DMemory_574 : _GEN_1690; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1692 = 10'h23f == EXMEMALUOut[9:0] ? DMemory_575 : _GEN_1691; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1693 = 10'h240 == EXMEMALUOut[9:0] ? DMemory_576 : _GEN_1692; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1694 = 10'h241 == EXMEMALUOut[9:0] ? DMemory_577 : _GEN_1693; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1695 = 10'h242 == EXMEMALUOut[9:0] ? DMemory_578 : _GEN_1694; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1696 = 10'h243 == EXMEMALUOut[9:0] ? DMemory_579 : _GEN_1695; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1697 = 10'h244 == EXMEMALUOut[9:0] ? DMemory_580 : _GEN_1696; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1698 = 10'h245 == EXMEMALUOut[9:0] ? DMemory_581 : _GEN_1697; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1699 = 10'h246 == EXMEMALUOut[9:0] ? DMemory_582 : _GEN_1698; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1700 = 10'h247 == EXMEMALUOut[9:0] ? DMemory_583 : _GEN_1699; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1701 = 10'h248 == EXMEMALUOut[9:0] ? DMemory_584 : _GEN_1700; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1702 = 10'h249 == EXMEMALUOut[9:0] ? DMemory_585 : _GEN_1701; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1703 = 10'h24a == EXMEMALUOut[9:0] ? DMemory_586 : _GEN_1702; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1704 = 10'h24b == EXMEMALUOut[9:0] ? DMemory_587 : _GEN_1703; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1705 = 10'h24c == EXMEMALUOut[9:0] ? DMemory_588 : _GEN_1704; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1706 = 10'h24d == EXMEMALUOut[9:0] ? DMemory_589 : _GEN_1705; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1707 = 10'h24e == EXMEMALUOut[9:0] ? DMemory_590 : _GEN_1706; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1708 = 10'h24f == EXMEMALUOut[9:0] ? DMemory_591 : _GEN_1707; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1709 = 10'h250 == EXMEMALUOut[9:0] ? DMemory_592 : _GEN_1708; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1710 = 10'h251 == EXMEMALUOut[9:0] ? DMemory_593 : _GEN_1709; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1711 = 10'h252 == EXMEMALUOut[9:0] ? DMemory_594 : _GEN_1710; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1712 = 10'h253 == EXMEMALUOut[9:0] ? DMemory_595 : _GEN_1711; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1713 = 10'h254 == EXMEMALUOut[9:0] ? DMemory_596 : _GEN_1712; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1714 = 10'h255 == EXMEMALUOut[9:0] ? DMemory_597 : _GEN_1713; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1715 = 10'h256 == EXMEMALUOut[9:0] ? DMemory_598 : _GEN_1714; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1716 = 10'h257 == EXMEMALUOut[9:0] ? DMemory_599 : _GEN_1715; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1717 = 10'h258 == EXMEMALUOut[9:0] ? DMemory_600 : _GEN_1716; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1718 = 10'h259 == EXMEMALUOut[9:0] ? DMemory_601 : _GEN_1717; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1719 = 10'h25a == EXMEMALUOut[9:0] ? DMemory_602 : _GEN_1718; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1720 = 10'h25b == EXMEMALUOut[9:0] ? DMemory_603 : _GEN_1719; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1721 = 10'h25c == EXMEMALUOut[9:0] ? DMemory_604 : _GEN_1720; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1722 = 10'h25d == EXMEMALUOut[9:0] ? DMemory_605 : _GEN_1721; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1723 = 10'h25e == EXMEMALUOut[9:0] ? DMemory_606 : _GEN_1722; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1724 = 10'h25f == EXMEMALUOut[9:0] ? DMemory_607 : _GEN_1723; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1725 = 10'h260 == EXMEMALUOut[9:0] ? DMemory_608 : _GEN_1724; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1726 = 10'h261 == EXMEMALUOut[9:0] ? DMemory_609 : _GEN_1725; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1727 = 10'h262 == EXMEMALUOut[9:0] ? DMemory_610 : _GEN_1726; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1728 = 10'h263 == EXMEMALUOut[9:0] ? DMemory_611 : _GEN_1727; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1729 = 10'h264 == EXMEMALUOut[9:0] ? DMemory_612 : _GEN_1728; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1730 = 10'h265 == EXMEMALUOut[9:0] ? DMemory_613 : _GEN_1729; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1731 = 10'h266 == EXMEMALUOut[9:0] ? DMemory_614 : _GEN_1730; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1732 = 10'h267 == EXMEMALUOut[9:0] ? DMemory_615 : _GEN_1731; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1733 = 10'h268 == EXMEMALUOut[9:0] ? DMemory_616 : _GEN_1732; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1734 = 10'h269 == EXMEMALUOut[9:0] ? DMemory_617 : _GEN_1733; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1735 = 10'h26a == EXMEMALUOut[9:0] ? DMemory_618 : _GEN_1734; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1736 = 10'h26b == EXMEMALUOut[9:0] ? DMemory_619 : _GEN_1735; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1737 = 10'h26c == EXMEMALUOut[9:0] ? DMemory_620 : _GEN_1736; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1738 = 10'h26d == EXMEMALUOut[9:0] ? DMemory_621 : _GEN_1737; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1739 = 10'h26e == EXMEMALUOut[9:0] ? DMemory_622 : _GEN_1738; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1740 = 10'h26f == EXMEMALUOut[9:0] ? DMemory_623 : _GEN_1739; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1741 = 10'h270 == EXMEMALUOut[9:0] ? DMemory_624 : _GEN_1740; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1742 = 10'h271 == EXMEMALUOut[9:0] ? DMemory_625 : _GEN_1741; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1743 = 10'h272 == EXMEMALUOut[9:0] ? DMemory_626 : _GEN_1742; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1744 = 10'h273 == EXMEMALUOut[9:0] ? DMemory_627 : _GEN_1743; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1745 = 10'h274 == EXMEMALUOut[9:0] ? DMemory_628 : _GEN_1744; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1746 = 10'h275 == EXMEMALUOut[9:0] ? DMemory_629 : _GEN_1745; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1747 = 10'h276 == EXMEMALUOut[9:0] ? DMemory_630 : _GEN_1746; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1748 = 10'h277 == EXMEMALUOut[9:0] ? DMemory_631 : _GEN_1747; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1749 = 10'h278 == EXMEMALUOut[9:0] ? DMemory_632 : _GEN_1748; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1750 = 10'h279 == EXMEMALUOut[9:0] ? DMemory_633 : _GEN_1749; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1751 = 10'h27a == EXMEMALUOut[9:0] ? DMemory_634 : _GEN_1750; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1752 = 10'h27b == EXMEMALUOut[9:0] ? DMemory_635 : _GEN_1751; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1753 = 10'h27c == EXMEMALUOut[9:0] ? DMemory_636 : _GEN_1752; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1754 = 10'h27d == EXMEMALUOut[9:0] ? DMemory_637 : _GEN_1753; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1755 = 10'h27e == EXMEMALUOut[9:0] ? DMemory_638 : _GEN_1754; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1756 = 10'h27f == EXMEMALUOut[9:0] ? DMemory_639 : _GEN_1755; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1757 = 10'h280 == EXMEMALUOut[9:0] ? DMemory_640 : _GEN_1756; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1758 = 10'h281 == EXMEMALUOut[9:0] ? DMemory_641 : _GEN_1757; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1759 = 10'h282 == EXMEMALUOut[9:0] ? DMemory_642 : _GEN_1758; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1760 = 10'h283 == EXMEMALUOut[9:0] ? DMemory_643 : _GEN_1759; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1761 = 10'h284 == EXMEMALUOut[9:0] ? DMemory_644 : _GEN_1760; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1762 = 10'h285 == EXMEMALUOut[9:0] ? DMemory_645 : _GEN_1761; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1763 = 10'h286 == EXMEMALUOut[9:0] ? DMemory_646 : _GEN_1762; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1764 = 10'h287 == EXMEMALUOut[9:0] ? DMemory_647 : _GEN_1763; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1765 = 10'h288 == EXMEMALUOut[9:0] ? DMemory_648 : _GEN_1764; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1766 = 10'h289 == EXMEMALUOut[9:0] ? DMemory_649 : _GEN_1765; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1767 = 10'h28a == EXMEMALUOut[9:0] ? DMemory_650 : _GEN_1766; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1768 = 10'h28b == EXMEMALUOut[9:0] ? DMemory_651 : _GEN_1767; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1769 = 10'h28c == EXMEMALUOut[9:0] ? DMemory_652 : _GEN_1768; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1770 = 10'h28d == EXMEMALUOut[9:0] ? DMemory_653 : _GEN_1769; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1771 = 10'h28e == EXMEMALUOut[9:0] ? DMemory_654 : _GEN_1770; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1772 = 10'h28f == EXMEMALUOut[9:0] ? DMemory_655 : _GEN_1771; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1773 = 10'h290 == EXMEMALUOut[9:0] ? DMemory_656 : _GEN_1772; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1774 = 10'h291 == EXMEMALUOut[9:0] ? DMemory_657 : _GEN_1773; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1775 = 10'h292 == EXMEMALUOut[9:0] ? DMemory_658 : _GEN_1774; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1776 = 10'h293 == EXMEMALUOut[9:0] ? DMemory_659 : _GEN_1775; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1777 = 10'h294 == EXMEMALUOut[9:0] ? DMemory_660 : _GEN_1776; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1778 = 10'h295 == EXMEMALUOut[9:0] ? DMemory_661 : _GEN_1777; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1779 = 10'h296 == EXMEMALUOut[9:0] ? DMemory_662 : _GEN_1778; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1780 = 10'h297 == EXMEMALUOut[9:0] ? DMemory_663 : _GEN_1779; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1781 = 10'h298 == EXMEMALUOut[9:0] ? DMemory_664 : _GEN_1780; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1782 = 10'h299 == EXMEMALUOut[9:0] ? DMemory_665 : _GEN_1781; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1783 = 10'h29a == EXMEMALUOut[9:0] ? DMemory_666 : _GEN_1782; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1784 = 10'h29b == EXMEMALUOut[9:0] ? DMemory_667 : _GEN_1783; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1785 = 10'h29c == EXMEMALUOut[9:0] ? DMemory_668 : _GEN_1784; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1786 = 10'h29d == EXMEMALUOut[9:0] ? DMemory_669 : _GEN_1785; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1787 = 10'h29e == EXMEMALUOut[9:0] ? DMemory_670 : _GEN_1786; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1788 = 10'h29f == EXMEMALUOut[9:0] ? DMemory_671 : _GEN_1787; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1789 = 10'h2a0 == EXMEMALUOut[9:0] ? DMemory_672 : _GEN_1788; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1790 = 10'h2a1 == EXMEMALUOut[9:0] ? DMemory_673 : _GEN_1789; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1791 = 10'h2a2 == EXMEMALUOut[9:0] ? DMemory_674 : _GEN_1790; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1792 = 10'h2a3 == EXMEMALUOut[9:0] ? DMemory_675 : _GEN_1791; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1793 = 10'h2a4 == EXMEMALUOut[9:0] ? DMemory_676 : _GEN_1792; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1794 = 10'h2a5 == EXMEMALUOut[9:0] ? DMemory_677 : _GEN_1793; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1795 = 10'h2a6 == EXMEMALUOut[9:0] ? DMemory_678 : _GEN_1794; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1796 = 10'h2a7 == EXMEMALUOut[9:0] ? DMemory_679 : _GEN_1795; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1797 = 10'h2a8 == EXMEMALUOut[9:0] ? DMemory_680 : _GEN_1796; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1798 = 10'h2a9 == EXMEMALUOut[9:0] ? DMemory_681 : _GEN_1797; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1799 = 10'h2aa == EXMEMALUOut[9:0] ? DMemory_682 : _GEN_1798; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1800 = 10'h2ab == EXMEMALUOut[9:0] ? DMemory_683 : _GEN_1799; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1801 = 10'h2ac == EXMEMALUOut[9:0] ? DMemory_684 : _GEN_1800; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1802 = 10'h2ad == EXMEMALUOut[9:0] ? DMemory_685 : _GEN_1801; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1803 = 10'h2ae == EXMEMALUOut[9:0] ? DMemory_686 : _GEN_1802; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1804 = 10'h2af == EXMEMALUOut[9:0] ? DMemory_687 : _GEN_1803; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1805 = 10'h2b0 == EXMEMALUOut[9:0] ? DMemory_688 : _GEN_1804; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1806 = 10'h2b1 == EXMEMALUOut[9:0] ? DMemory_689 : _GEN_1805; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1807 = 10'h2b2 == EXMEMALUOut[9:0] ? DMemory_690 : _GEN_1806; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1808 = 10'h2b3 == EXMEMALUOut[9:0] ? DMemory_691 : _GEN_1807; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1809 = 10'h2b4 == EXMEMALUOut[9:0] ? DMemory_692 : _GEN_1808; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1810 = 10'h2b5 == EXMEMALUOut[9:0] ? DMemory_693 : _GEN_1809; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1811 = 10'h2b6 == EXMEMALUOut[9:0] ? DMemory_694 : _GEN_1810; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1812 = 10'h2b7 == EXMEMALUOut[9:0] ? DMemory_695 : _GEN_1811; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1813 = 10'h2b8 == EXMEMALUOut[9:0] ? DMemory_696 : _GEN_1812; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1814 = 10'h2b9 == EXMEMALUOut[9:0] ? DMemory_697 : _GEN_1813; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1815 = 10'h2ba == EXMEMALUOut[9:0] ? DMemory_698 : _GEN_1814; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1816 = 10'h2bb == EXMEMALUOut[9:0] ? DMemory_699 : _GEN_1815; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1817 = 10'h2bc == EXMEMALUOut[9:0] ? DMemory_700 : _GEN_1816; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1818 = 10'h2bd == EXMEMALUOut[9:0] ? DMemory_701 : _GEN_1817; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1819 = 10'h2be == EXMEMALUOut[9:0] ? DMemory_702 : _GEN_1818; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1820 = 10'h2bf == EXMEMALUOut[9:0] ? DMemory_703 : _GEN_1819; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1821 = 10'h2c0 == EXMEMALUOut[9:0] ? DMemory_704 : _GEN_1820; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1822 = 10'h2c1 == EXMEMALUOut[9:0] ? DMemory_705 : _GEN_1821; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1823 = 10'h2c2 == EXMEMALUOut[9:0] ? DMemory_706 : _GEN_1822; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1824 = 10'h2c3 == EXMEMALUOut[9:0] ? DMemory_707 : _GEN_1823; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1825 = 10'h2c4 == EXMEMALUOut[9:0] ? DMemory_708 : _GEN_1824; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1826 = 10'h2c5 == EXMEMALUOut[9:0] ? DMemory_709 : _GEN_1825; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1827 = 10'h2c6 == EXMEMALUOut[9:0] ? DMemory_710 : _GEN_1826; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1828 = 10'h2c7 == EXMEMALUOut[9:0] ? DMemory_711 : _GEN_1827; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1829 = 10'h2c8 == EXMEMALUOut[9:0] ? DMemory_712 : _GEN_1828; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1830 = 10'h2c9 == EXMEMALUOut[9:0] ? DMemory_713 : _GEN_1829; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1831 = 10'h2ca == EXMEMALUOut[9:0] ? DMemory_714 : _GEN_1830; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1832 = 10'h2cb == EXMEMALUOut[9:0] ? DMemory_715 : _GEN_1831; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1833 = 10'h2cc == EXMEMALUOut[9:0] ? DMemory_716 : _GEN_1832; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1834 = 10'h2cd == EXMEMALUOut[9:0] ? DMemory_717 : _GEN_1833; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1835 = 10'h2ce == EXMEMALUOut[9:0] ? DMemory_718 : _GEN_1834; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1836 = 10'h2cf == EXMEMALUOut[9:0] ? DMemory_719 : _GEN_1835; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1837 = 10'h2d0 == EXMEMALUOut[9:0] ? DMemory_720 : _GEN_1836; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1838 = 10'h2d1 == EXMEMALUOut[9:0] ? DMemory_721 : _GEN_1837; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1839 = 10'h2d2 == EXMEMALUOut[9:0] ? DMemory_722 : _GEN_1838; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1840 = 10'h2d3 == EXMEMALUOut[9:0] ? DMemory_723 : _GEN_1839; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1841 = 10'h2d4 == EXMEMALUOut[9:0] ? DMemory_724 : _GEN_1840; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1842 = 10'h2d5 == EXMEMALUOut[9:0] ? DMemory_725 : _GEN_1841; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1843 = 10'h2d6 == EXMEMALUOut[9:0] ? DMemory_726 : _GEN_1842; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1844 = 10'h2d7 == EXMEMALUOut[9:0] ? DMemory_727 : _GEN_1843; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1845 = 10'h2d8 == EXMEMALUOut[9:0] ? DMemory_728 : _GEN_1844; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1846 = 10'h2d9 == EXMEMALUOut[9:0] ? DMemory_729 : _GEN_1845; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1847 = 10'h2da == EXMEMALUOut[9:0] ? DMemory_730 : _GEN_1846; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1848 = 10'h2db == EXMEMALUOut[9:0] ? DMemory_731 : _GEN_1847; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1849 = 10'h2dc == EXMEMALUOut[9:0] ? DMemory_732 : _GEN_1848; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1850 = 10'h2dd == EXMEMALUOut[9:0] ? DMemory_733 : _GEN_1849; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1851 = 10'h2de == EXMEMALUOut[9:0] ? DMemory_734 : _GEN_1850; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1852 = 10'h2df == EXMEMALUOut[9:0] ? DMemory_735 : _GEN_1851; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1853 = 10'h2e0 == EXMEMALUOut[9:0] ? DMemory_736 : _GEN_1852; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1854 = 10'h2e1 == EXMEMALUOut[9:0] ? DMemory_737 : _GEN_1853; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1855 = 10'h2e2 == EXMEMALUOut[9:0] ? DMemory_738 : _GEN_1854; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1856 = 10'h2e3 == EXMEMALUOut[9:0] ? DMemory_739 : _GEN_1855; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1857 = 10'h2e4 == EXMEMALUOut[9:0] ? DMemory_740 : _GEN_1856; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1858 = 10'h2e5 == EXMEMALUOut[9:0] ? DMemory_741 : _GEN_1857; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1859 = 10'h2e6 == EXMEMALUOut[9:0] ? DMemory_742 : _GEN_1858; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1860 = 10'h2e7 == EXMEMALUOut[9:0] ? DMemory_743 : _GEN_1859; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1861 = 10'h2e8 == EXMEMALUOut[9:0] ? DMemory_744 : _GEN_1860; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1862 = 10'h2e9 == EXMEMALUOut[9:0] ? DMemory_745 : _GEN_1861; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1863 = 10'h2ea == EXMEMALUOut[9:0] ? DMemory_746 : _GEN_1862; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1864 = 10'h2eb == EXMEMALUOut[9:0] ? DMemory_747 : _GEN_1863; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1865 = 10'h2ec == EXMEMALUOut[9:0] ? DMemory_748 : _GEN_1864; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1866 = 10'h2ed == EXMEMALUOut[9:0] ? DMemory_749 : _GEN_1865; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1867 = 10'h2ee == EXMEMALUOut[9:0] ? DMemory_750 : _GEN_1866; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1868 = 10'h2ef == EXMEMALUOut[9:0] ? DMemory_751 : _GEN_1867; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1869 = 10'h2f0 == EXMEMALUOut[9:0] ? DMemory_752 : _GEN_1868; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1870 = 10'h2f1 == EXMEMALUOut[9:0] ? DMemory_753 : _GEN_1869; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1871 = 10'h2f2 == EXMEMALUOut[9:0] ? DMemory_754 : _GEN_1870; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1872 = 10'h2f3 == EXMEMALUOut[9:0] ? DMemory_755 : _GEN_1871; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1873 = 10'h2f4 == EXMEMALUOut[9:0] ? DMemory_756 : _GEN_1872; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1874 = 10'h2f5 == EXMEMALUOut[9:0] ? DMemory_757 : _GEN_1873; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1875 = 10'h2f6 == EXMEMALUOut[9:0] ? DMemory_758 : _GEN_1874; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1876 = 10'h2f7 == EXMEMALUOut[9:0] ? DMemory_759 : _GEN_1875; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1877 = 10'h2f8 == EXMEMALUOut[9:0] ? DMemory_760 : _GEN_1876; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1878 = 10'h2f9 == EXMEMALUOut[9:0] ? DMemory_761 : _GEN_1877; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1879 = 10'h2fa == EXMEMALUOut[9:0] ? DMemory_762 : _GEN_1878; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1880 = 10'h2fb == EXMEMALUOut[9:0] ? DMemory_763 : _GEN_1879; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1881 = 10'h2fc == EXMEMALUOut[9:0] ? DMemory_764 : _GEN_1880; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1882 = 10'h2fd == EXMEMALUOut[9:0] ? DMemory_765 : _GEN_1881; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1883 = 10'h2fe == EXMEMALUOut[9:0] ? DMemory_766 : _GEN_1882; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1884 = 10'h2ff == EXMEMALUOut[9:0] ? DMemory_767 : _GEN_1883; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1885 = 10'h300 == EXMEMALUOut[9:0] ? DMemory_768 : _GEN_1884; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1886 = 10'h301 == EXMEMALUOut[9:0] ? DMemory_769 : _GEN_1885; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1887 = 10'h302 == EXMEMALUOut[9:0] ? DMemory_770 : _GEN_1886; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1888 = 10'h303 == EXMEMALUOut[9:0] ? DMemory_771 : _GEN_1887; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1889 = 10'h304 == EXMEMALUOut[9:0] ? DMemory_772 : _GEN_1888; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1890 = 10'h305 == EXMEMALUOut[9:0] ? DMemory_773 : _GEN_1889; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1891 = 10'h306 == EXMEMALUOut[9:0] ? DMemory_774 : _GEN_1890; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1892 = 10'h307 == EXMEMALUOut[9:0] ? DMemory_775 : _GEN_1891; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1893 = 10'h308 == EXMEMALUOut[9:0] ? DMemory_776 : _GEN_1892; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1894 = 10'h309 == EXMEMALUOut[9:0] ? DMemory_777 : _GEN_1893; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1895 = 10'h30a == EXMEMALUOut[9:0] ? DMemory_778 : _GEN_1894; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1896 = 10'h30b == EXMEMALUOut[9:0] ? DMemory_779 : _GEN_1895; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1897 = 10'h30c == EXMEMALUOut[9:0] ? DMemory_780 : _GEN_1896; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1898 = 10'h30d == EXMEMALUOut[9:0] ? DMemory_781 : _GEN_1897; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1899 = 10'h30e == EXMEMALUOut[9:0] ? DMemory_782 : _GEN_1898; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1900 = 10'h30f == EXMEMALUOut[9:0] ? DMemory_783 : _GEN_1899; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1901 = 10'h310 == EXMEMALUOut[9:0] ? DMemory_784 : _GEN_1900; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1902 = 10'h311 == EXMEMALUOut[9:0] ? DMemory_785 : _GEN_1901; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1903 = 10'h312 == EXMEMALUOut[9:0] ? DMemory_786 : _GEN_1902; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1904 = 10'h313 == EXMEMALUOut[9:0] ? DMemory_787 : _GEN_1903; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1905 = 10'h314 == EXMEMALUOut[9:0] ? DMemory_788 : _GEN_1904; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1906 = 10'h315 == EXMEMALUOut[9:0] ? DMemory_789 : _GEN_1905; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1907 = 10'h316 == EXMEMALUOut[9:0] ? DMemory_790 : _GEN_1906; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1908 = 10'h317 == EXMEMALUOut[9:0] ? DMemory_791 : _GEN_1907; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1909 = 10'h318 == EXMEMALUOut[9:0] ? DMemory_792 : _GEN_1908; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1910 = 10'h319 == EXMEMALUOut[9:0] ? DMemory_793 : _GEN_1909; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1911 = 10'h31a == EXMEMALUOut[9:0] ? DMemory_794 : _GEN_1910; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1912 = 10'h31b == EXMEMALUOut[9:0] ? DMemory_795 : _GEN_1911; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1913 = 10'h31c == EXMEMALUOut[9:0] ? DMemory_796 : _GEN_1912; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1914 = 10'h31d == EXMEMALUOut[9:0] ? DMemory_797 : _GEN_1913; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1915 = 10'h31e == EXMEMALUOut[9:0] ? DMemory_798 : _GEN_1914; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1916 = 10'h31f == EXMEMALUOut[9:0] ? DMemory_799 : _GEN_1915; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1917 = 10'h320 == EXMEMALUOut[9:0] ? DMemory_800 : _GEN_1916; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1918 = 10'h321 == EXMEMALUOut[9:0] ? DMemory_801 : _GEN_1917; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1919 = 10'h322 == EXMEMALUOut[9:0] ? DMemory_802 : _GEN_1918; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1920 = 10'h323 == EXMEMALUOut[9:0] ? DMemory_803 : _GEN_1919; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1921 = 10'h324 == EXMEMALUOut[9:0] ? DMemory_804 : _GEN_1920; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1922 = 10'h325 == EXMEMALUOut[9:0] ? DMemory_805 : _GEN_1921; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1923 = 10'h326 == EXMEMALUOut[9:0] ? DMemory_806 : _GEN_1922; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1924 = 10'h327 == EXMEMALUOut[9:0] ? DMemory_807 : _GEN_1923; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1925 = 10'h328 == EXMEMALUOut[9:0] ? DMemory_808 : _GEN_1924; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1926 = 10'h329 == EXMEMALUOut[9:0] ? DMemory_809 : _GEN_1925; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1927 = 10'h32a == EXMEMALUOut[9:0] ? DMemory_810 : _GEN_1926; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1928 = 10'h32b == EXMEMALUOut[9:0] ? DMemory_811 : _GEN_1927; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1929 = 10'h32c == EXMEMALUOut[9:0] ? DMemory_812 : _GEN_1928; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1930 = 10'h32d == EXMEMALUOut[9:0] ? DMemory_813 : _GEN_1929; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1931 = 10'h32e == EXMEMALUOut[9:0] ? DMemory_814 : _GEN_1930; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1932 = 10'h32f == EXMEMALUOut[9:0] ? DMemory_815 : _GEN_1931; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1933 = 10'h330 == EXMEMALUOut[9:0] ? DMemory_816 : _GEN_1932; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1934 = 10'h331 == EXMEMALUOut[9:0] ? DMemory_817 : _GEN_1933; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1935 = 10'h332 == EXMEMALUOut[9:0] ? DMemory_818 : _GEN_1934; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1936 = 10'h333 == EXMEMALUOut[9:0] ? DMemory_819 : _GEN_1935; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1937 = 10'h334 == EXMEMALUOut[9:0] ? DMemory_820 : _GEN_1936; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1938 = 10'h335 == EXMEMALUOut[9:0] ? DMemory_821 : _GEN_1937; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1939 = 10'h336 == EXMEMALUOut[9:0] ? DMemory_822 : _GEN_1938; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1940 = 10'h337 == EXMEMALUOut[9:0] ? DMemory_823 : _GEN_1939; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1941 = 10'h338 == EXMEMALUOut[9:0] ? DMemory_824 : _GEN_1940; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1942 = 10'h339 == EXMEMALUOut[9:0] ? DMemory_825 : _GEN_1941; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1943 = 10'h33a == EXMEMALUOut[9:0] ? DMemory_826 : _GEN_1942; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1944 = 10'h33b == EXMEMALUOut[9:0] ? DMemory_827 : _GEN_1943; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1945 = 10'h33c == EXMEMALUOut[9:0] ? DMemory_828 : _GEN_1944; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1946 = 10'h33d == EXMEMALUOut[9:0] ? DMemory_829 : _GEN_1945; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1947 = 10'h33e == EXMEMALUOut[9:0] ? DMemory_830 : _GEN_1946; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1948 = 10'h33f == EXMEMALUOut[9:0] ? DMemory_831 : _GEN_1947; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1949 = 10'h340 == EXMEMALUOut[9:0] ? DMemory_832 : _GEN_1948; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1950 = 10'h341 == EXMEMALUOut[9:0] ? DMemory_833 : _GEN_1949; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1951 = 10'h342 == EXMEMALUOut[9:0] ? DMemory_834 : _GEN_1950; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1952 = 10'h343 == EXMEMALUOut[9:0] ? DMemory_835 : _GEN_1951; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1953 = 10'h344 == EXMEMALUOut[9:0] ? DMemory_836 : _GEN_1952; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1954 = 10'h345 == EXMEMALUOut[9:0] ? DMemory_837 : _GEN_1953; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1955 = 10'h346 == EXMEMALUOut[9:0] ? DMemory_838 : _GEN_1954; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1956 = 10'h347 == EXMEMALUOut[9:0] ? DMemory_839 : _GEN_1955; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1957 = 10'h348 == EXMEMALUOut[9:0] ? DMemory_840 : _GEN_1956; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1958 = 10'h349 == EXMEMALUOut[9:0] ? DMemory_841 : _GEN_1957; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1959 = 10'h34a == EXMEMALUOut[9:0] ? DMemory_842 : _GEN_1958; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1960 = 10'h34b == EXMEMALUOut[9:0] ? DMemory_843 : _GEN_1959; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1961 = 10'h34c == EXMEMALUOut[9:0] ? DMemory_844 : _GEN_1960; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1962 = 10'h34d == EXMEMALUOut[9:0] ? DMemory_845 : _GEN_1961; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1963 = 10'h34e == EXMEMALUOut[9:0] ? DMemory_846 : _GEN_1962; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1964 = 10'h34f == EXMEMALUOut[9:0] ? DMemory_847 : _GEN_1963; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1965 = 10'h350 == EXMEMALUOut[9:0] ? DMemory_848 : _GEN_1964; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1966 = 10'h351 == EXMEMALUOut[9:0] ? DMemory_849 : _GEN_1965; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1967 = 10'h352 == EXMEMALUOut[9:0] ? DMemory_850 : _GEN_1966; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1968 = 10'h353 == EXMEMALUOut[9:0] ? DMemory_851 : _GEN_1967; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1969 = 10'h354 == EXMEMALUOut[9:0] ? DMemory_852 : _GEN_1968; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1970 = 10'h355 == EXMEMALUOut[9:0] ? DMemory_853 : _GEN_1969; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1971 = 10'h356 == EXMEMALUOut[9:0] ? DMemory_854 : _GEN_1970; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1972 = 10'h357 == EXMEMALUOut[9:0] ? DMemory_855 : _GEN_1971; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1973 = 10'h358 == EXMEMALUOut[9:0] ? DMemory_856 : _GEN_1972; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1974 = 10'h359 == EXMEMALUOut[9:0] ? DMemory_857 : _GEN_1973; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1975 = 10'h35a == EXMEMALUOut[9:0] ? DMemory_858 : _GEN_1974; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1976 = 10'h35b == EXMEMALUOut[9:0] ? DMemory_859 : _GEN_1975; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1977 = 10'h35c == EXMEMALUOut[9:0] ? DMemory_860 : _GEN_1976; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1978 = 10'h35d == EXMEMALUOut[9:0] ? DMemory_861 : _GEN_1977; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1979 = 10'h35e == EXMEMALUOut[9:0] ? DMemory_862 : _GEN_1978; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1980 = 10'h35f == EXMEMALUOut[9:0] ? DMemory_863 : _GEN_1979; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1981 = 10'h360 == EXMEMALUOut[9:0] ? DMemory_864 : _GEN_1980; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1982 = 10'h361 == EXMEMALUOut[9:0] ? DMemory_865 : _GEN_1981; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1983 = 10'h362 == EXMEMALUOut[9:0] ? DMemory_866 : _GEN_1982; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1984 = 10'h363 == EXMEMALUOut[9:0] ? DMemory_867 : _GEN_1983; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1985 = 10'h364 == EXMEMALUOut[9:0] ? DMemory_868 : _GEN_1984; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1986 = 10'h365 == EXMEMALUOut[9:0] ? DMemory_869 : _GEN_1985; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1987 = 10'h366 == EXMEMALUOut[9:0] ? DMemory_870 : _GEN_1986; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1988 = 10'h367 == EXMEMALUOut[9:0] ? DMemory_871 : _GEN_1987; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1989 = 10'h368 == EXMEMALUOut[9:0] ? DMemory_872 : _GEN_1988; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1990 = 10'h369 == EXMEMALUOut[9:0] ? DMemory_873 : _GEN_1989; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1991 = 10'h36a == EXMEMALUOut[9:0] ? DMemory_874 : _GEN_1990; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1992 = 10'h36b == EXMEMALUOut[9:0] ? DMemory_875 : _GEN_1991; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1993 = 10'h36c == EXMEMALUOut[9:0] ? DMemory_876 : _GEN_1992; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1994 = 10'h36d == EXMEMALUOut[9:0] ? DMemory_877 : _GEN_1993; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1995 = 10'h36e == EXMEMALUOut[9:0] ? DMemory_878 : _GEN_1994; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1996 = 10'h36f == EXMEMALUOut[9:0] ? DMemory_879 : _GEN_1995; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1997 = 10'h370 == EXMEMALUOut[9:0] ? DMemory_880 : _GEN_1996; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1998 = 10'h371 == EXMEMALUOut[9:0] ? DMemory_881 : _GEN_1997; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_1999 = 10'h372 == EXMEMALUOut[9:0] ? DMemory_882 : _GEN_1998; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2000 = 10'h373 == EXMEMALUOut[9:0] ? DMemory_883 : _GEN_1999; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2001 = 10'h374 == EXMEMALUOut[9:0] ? DMemory_884 : _GEN_2000; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2002 = 10'h375 == EXMEMALUOut[9:0] ? DMemory_885 : _GEN_2001; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2003 = 10'h376 == EXMEMALUOut[9:0] ? DMemory_886 : _GEN_2002; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2004 = 10'h377 == EXMEMALUOut[9:0] ? DMemory_887 : _GEN_2003; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2005 = 10'h378 == EXMEMALUOut[9:0] ? DMemory_888 : _GEN_2004; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2006 = 10'h379 == EXMEMALUOut[9:0] ? DMemory_889 : _GEN_2005; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2007 = 10'h37a == EXMEMALUOut[9:0] ? DMemory_890 : _GEN_2006; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2008 = 10'h37b == EXMEMALUOut[9:0] ? DMemory_891 : _GEN_2007; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2009 = 10'h37c == EXMEMALUOut[9:0] ? DMemory_892 : _GEN_2008; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2010 = 10'h37d == EXMEMALUOut[9:0] ? DMemory_893 : _GEN_2009; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2011 = 10'h37e == EXMEMALUOut[9:0] ? DMemory_894 : _GEN_2010; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2012 = 10'h37f == EXMEMALUOut[9:0] ? DMemory_895 : _GEN_2011; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2013 = 10'h380 == EXMEMALUOut[9:0] ? DMemory_896 : _GEN_2012; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2014 = 10'h381 == EXMEMALUOut[9:0] ? DMemory_897 : _GEN_2013; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2015 = 10'h382 == EXMEMALUOut[9:0] ? DMemory_898 : _GEN_2014; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2016 = 10'h383 == EXMEMALUOut[9:0] ? DMemory_899 : _GEN_2015; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2017 = 10'h384 == EXMEMALUOut[9:0] ? DMemory_900 : _GEN_2016; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2018 = 10'h385 == EXMEMALUOut[9:0] ? DMemory_901 : _GEN_2017; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2019 = 10'h386 == EXMEMALUOut[9:0] ? DMemory_902 : _GEN_2018; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2020 = 10'h387 == EXMEMALUOut[9:0] ? DMemory_903 : _GEN_2019; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2021 = 10'h388 == EXMEMALUOut[9:0] ? DMemory_904 : _GEN_2020; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2022 = 10'h389 == EXMEMALUOut[9:0] ? DMemory_905 : _GEN_2021; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2023 = 10'h38a == EXMEMALUOut[9:0] ? DMemory_906 : _GEN_2022; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2024 = 10'h38b == EXMEMALUOut[9:0] ? DMemory_907 : _GEN_2023; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2025 = 10'h38c == EXMEMALUOut[9:0] ? DMemory_908 : _GEN_2024; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2026 = 10'h38d == EXMEMALUOut[9:0] ? DMemory_909 : _GEN_2025; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2027 = 10'h38e == EXMEMALUOut[9:0] ? DMemory_910 : _GEN_2026; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2028 = 10'h38f == EXMEMALUOut[9:0] ? DMemory_911 : _GEN_2027; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2029 = 10'h390 == EXMEMALUOut[9:0] ? DMemory_912 : _GEN_2028; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2030 = 10'h391 == EXMEMALUOut[9:0] ? DMemory_913 : _GEN_2029; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2031 = 10'h392 == EXMEMALUOut[9:0] ? DMemory_914 : _GEN_2030; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2032 = 10'h393 == EXMEMALUOut[9:0] ? DMemory_915 : _GEN_2031; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2033 = 10'h394 == EXMEMALUOut[9:0] ? DMemory_916 : _GEN_2032; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2034 = 10'h395 == EXMEMALUOut[9:0] ? DMemory_917 : _GEN_2033; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2035 = 10'h396 == EXMEMALUOut[9:0] ? DMemory_918 : _GEN_2034; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2036 = 10'h397 == EXMEMALUOut[9:0] ? DMemory_919 : _GEN_2035; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2037 = 10'h398 == EXMEMALUOut[9:0] ? DMemory_920 : _GEN_2036; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2038 = 10'h399 == EXMEMALUOut[9:0] ? DMemory_921 : _GEN_2037; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2039 = 10'h39a == EXMEMALUOut[9:0] ? DMemory_922 : _GEN_2038; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2040 = 10'h39b == EXMEMALUOut[9:0] ? DMemory_923 : _GEN_2039; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2041 = 10'h39c == EXMEMALUOut[9:0] ? DMemory_924 : _GEN_2040; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2042 = 10'h39d == EXMEMALUOut[9:0] ? DMemory_925 : _GEN_2041; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2043 = 10'h39e == EXMEMALUOut[9:0] ? DMemory_926 : _GEN_2042; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2044 = 10'h39f == EXMEMALUOut[9:0] ? DMemory_927 : _GEN_2043; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2045 = 10'h3a0 == EXMEMALUOut[9:0] ? DMemory_928 : _GEN_2044; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2046 = 10'h3a1 == EXMEMALUOut[9:0] ? DMemory_929 : _GEN_2045; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2047 = 10'h3a2 == EXMEMALUOut[9:0] ? DMemory_930 : _GEN_2046; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2048 = 10'h3a3 == EXMEMALUOut[9:0] ? DMemory_931 : _GEN_2047; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2049 = 10'h3a4 == EXMEMALUOut[9:0] ? DMemory_932 : _GEN_2048; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2050 = 10'h3a5 == EXMEMALUOut[9:0] ? DMemory_933 : _GEN_2049; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2051 = 10'h3a6 == EXMEMALUOut[9:0] ? DMemory_934 : _GEN_2050; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2052 = 10'h3a7 == EXMEMALUOut[9:0] ? DMemory_935 : _GEN_2051; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2053 = 10'h3a8 == EXMEMALUOut[9:0] ? DMemory_936 : _GEN_2052; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2054 = 10'h3a9 == EXMEMALUOut[9:0] ? DMemory_937 : _GEN_2053; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2055 = 10'h3aa == EXMEMALUOut[9:0] ? DMemory_938 : _GEN_2054; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2056 = 10'h3ab == EXMEMALUOut[9:0] ? DMemory_939 : _GEN_2055; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2057 = 10'h3ac == EXMEMALUOut[9:0] ? DMemory_940 : _GEN_2056; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2058 = 10'h3ad == EXMEMALUOut[9:0] ? DMemory_941 : _GEN_2057; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2059 = 10'h3ae == EXMEMALUOut[9:0] ? DMemory_942 : _GEN_2058; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2060 = 10'h3af == EXMEMALUOut[9:0] ? DMemory_943 : _GEN_2059; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2061 = 10'h3b0 == EXMEMALUOut[9:0] ? DMemory_944 : _GEN_2060; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2062 = 10'h3b1 == EXMEMALUOut[9:0] ? DMemory_945 : _GEN_2061; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2063 = 10'h3b2 == EXMEMALUOut[9:0] ? DMemory_946 : _GEN_2062; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2064 = 10'h3b3 == EXMEMALUOut[9:0] ? DMemory_947 : _GEN_2063; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2065 = 10'h3b4 == EXMEMALUOut[9:0] ? DMemory_948 : _GEN_2064; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2066 = 10'h3b5 == EXMEMALUOut[9:0] ? DMemory_949 : _GEN_2065; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2067 = 10'h3b6 == EXMEMALUOut[9:0] ? DMemory_950 : _GEN_2066; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2068 = 10'h3b7 == EXMEMALUOut[9:0] ? DMemory_951 : _GEN_2067; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2069 = 10'h3b8 == EXMEMALUOut[9:0] ? DMemory_952 : _GEN_2068; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2070 = 10'h3b9 == EXMEMALUOut[9:0] ? DMemory_953 : _GEN_2069; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2071 = 10'h3ba == EXMEMALUOut[9:0] ? DMemory_954 : _GEN_2070; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2072 = 10'h3bb == EXMEMALUOut[9:0] ? DMemory_955 : _GEN_2071; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2073 = 10'h3bc == EXMEMALUOut[9:0] ? DMemory_956 : _GEN_2072; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2074 = 10'h3bd == EXMEMALUOut[9:0] ? DMemory_957 : _GEN_2073; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2075 = 10'h3be == EXMEMALUOut[9:0] ? DMemory_958 : _GEN_2074; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2076 = 10'h3bf == EXMEMALUOut[9:0] ? DMemory_959 : _GEN_2075; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2077 = 10'h3c0 == EXMEMALUOut[9:0] ? DMemory_960 : _GEN_2076; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2078 = 10'h3c1 == EXMEMALUOut[9:0] ? DMemory_961 : _GEN_2077; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2079 = 10'h3c2 == EXMEMALUOut[9:0] ? DMemory_962 : _GEN_2078; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2080 = 10'h3c3 == EXMEMALUOut[9:0] ? DMemory_963 : _GEN_2079; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2081 = 10'h3c4 == EXMEMALUOut[9:0] ? DMemory_964 : _GEN_2080; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2082 = 10'h3c5 == EXMEMALUOut[9:0] ? DMemory_965 : _GEN_2081; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2083 = 10'h3c6 == EXMEMALUOut[9:0] ? DMemory_966 : _GEN_2082; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2084 = 10'h3c7 == EXMEMALUOut[9:0] ? DMemory_967 : _GEN_2083; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2085 = 10'h3c8 == EXMEMALUOut[9:0] ? DMemory_968 : _GEN_2084; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2086 = 10'h3c9 == EXMEMALUOut[9:0] ? DMemory_969 : _GEN_2085; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2087 = 10'h3ca == EXMEMALUOut[9:0] ? DMemory_970 : _GEN_2086; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2088 = 10'h3cb == EXMEMALUOut[9:0] ? DMemory_971 : _GEN_2087; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2089 = 10'h3cc == EXMEMALUOut[9:0] ? DMemory_972 : _GEN_2088; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2090 = 10'h3cd == EXMEMALUOut[9:0] ? DMemory_973 : _GEN_2089; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2091 = 10'h3ce == EXMEMALUOut[9:0] ? DMemory_974 : _GEN_2090; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2092 = 10'h3cf == EXMEMALUOut[9:0] ? DMemory_975 : _GEN_2091; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2093 = 10'h3d0 == EXMEMALUOut[9:0] ? DMemory_976 : _GEN_2092; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2094 = 10'h3d1 == EXMEMALUOut[9:0] ? DMemory_977 : _GEN_2093; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2095 = 10'h3d2 == EXMEMALUOut[9:0] ? DMemory_978 : _GEN_2094; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2096 = 10'h3d3 == EXMEMALUOut[9:0] ? DMemory_979 : _GEN_2095; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2097 = 10'h3d4 == EXMEMALUOut[9:0] ? DMemory_980 : _GEN_2096; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2098 = 10'h3d5 == EXMEMALUOut[9:0] ? DMemory_981 : _GEN_2097; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2099 = 10'h3d6 == EXMEMALUOut[9:0] ? DMemory_982 : _GEN_2098; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2100 = 10'h3d7 == EXMEMALUOut[9:0] ? DMemory_983 : _GEN_2099; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2101 = 10'h3d8 == EXMEMALUOut[9:0] ? DMemory_984 : _GEN_2100; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2102 = 10'h3d9 == EXMEMALUOut[9:0] ? DMemory_985 : _GEN_2101; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2103 = 10'h3da == EXMEMALUOut[9:0] ? DMemory_986 : _GEN_2102; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2104 = 10'h3db == EXMEMALUOut[9:0] ? DMemory_987 : _GEN_2103; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2105 = 10'h3dc == EXMEMALUOut[9:0] ? DMemory_988 : _GEN_2104; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2106 = 10'h3dd == EXMEMALUOut[9:0] ? DMemory_989 : _GEN_2105; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2107 = 10'h3de == EXMEMALUOut[9:0] ? DMemory_990 : _GEN_2106; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2108 = 10'h3df == EXMEMALUOut[9:0] ? DMemory_991 : _GEN_2107; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2109 = 10'h3e0 == EXMEMALUOut[9:0] ? DMemory_992 : _GEN_2108; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2110 = 10'h3e1 == EXMEMALUOut[9:0] ? DMemory_993 : _GEN_2109; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2111 = 10'h3e2 == EXMEMALUOut[9:0] ? DMemory_994 : _GEN_2110; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2112 = 10'h3e3 == EXMEMALUOut[9:0] ? DMemory_995 : _GEN_2111; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2113 = 10'h3e4 == EXMEMALUOut[9:0] ? DMemory_996 : _GEN_2112; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2114 = 10'h3e5 == EXMEMALUOut[9:0] ? DMemory_997 : _GEN_2113; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2115 = 10'h3e6 == EXMEMALUOut[9:0] ? DMemory_998 : _GEN_2114; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2116 = 10'h3e7 == EXMEMALUOut[9:0] ? DMemory_999 : _GEN_2115; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2117 = 10'h3e8 == EXMEMALUOut[9:0] ? DMemory_1000 : _GEN_2116; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2118 = 10'h3e9 == EXMEMALUOut[9:0] ? DMemory_1001 : _GEN_2117; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2119 = 10'h3ea == EXMEMALUOut[9:0] ? DMemory_1002 : _GEN_2118; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2120 = 10'h3eb == EXMEMALUOut[9:0] ? DMemory_1003 : _GEN_2119; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2121 = 10'h3ec == EXMEMALUOut[9:0] ? DMemory_1004 : _GEN_2120; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2122 = 10'h3ed == EXMEMALUOut[9:0] ? DMemory_1005 : _GEN_2121; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2123 = 10'h3ee == EXMEMALUOut[9:0] ? DMemory_1006 : _GEN_2122; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2124 = 10'h3ef == EXMEMALUOut[9:0] ? DMemory_1007 : _GEN_2123; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2125 = 10'h3f0 == EXMEMALUOut[9:0] ? DMemory_1008 : _GEN_2124; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2126 = 10'h3f1 == EXMEMALUOut[9:0] ? DMemory_1009 : _GEN_2125; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2127 = 10'h3f2 == EXMEMALUOut[9:0] ? DMemory_1010 : _GEN_2126; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2128 = 10'h3f3 == EXMEMALUOut[9:0] ? DMemory_1011 : _GEN_2127; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2129 = 10'h3f4 == EXMEMALUOut[9:0] ? DMemory_1012 : _GEN_2128; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2130 = 10'h3f5 == EXMEMALUOut[9:0] ? DMemory_1013 : _GEN_2129; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2131 = 10'h3f6 == EXMEMALUOut[9:0] ? DMemory_1014 : _GEN_2130; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2132 = 10'h3f7 == EXMEMALUOut[9:0] ? DMemory_1015 : _GEN_2131; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2133 = 10'h3f8 == EXMEMALUOut[9:0] ? DMemory_1016 : _GEN_2132; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2134 = 10'h3f9 == EXMEMALUOut[9:0] ? DMemory_1017 : _GEN_2133; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2135 = 10'h3fa == EXMEMALUOut[9:0] ? DMemory_1018 : _GEN_2134; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2136 = 10'h3fb == EXMEMALUOut[9:0] ? DMemory_1019 : _GEN_2135; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2137 = 10'h3fc == EXMEMALUOut[9:0] ? DMemory_1020 : _GEN_2136; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2138 = 10'h3fd == EXMEMALUOut[9:0] ? DMemory_1021 : _GEN_2137; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2139 = 10'h3fe == EXMEMALUOut[9:0] ? DMemory_1022 : _GEN_2138; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2140 = 10'h3ff == EXMEMALUOut[9:0] ? DMemory_1023 : _GEN_2139; // @[cpu.scala 199:{18,18}]
  wire [31:0] _GEN_2141 = 10'h0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_0; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2142 = 10'h1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2143 = 10'h2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_2; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2144 = 10'h3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_3; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2145 = 10'h4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_4; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2146 = 10'h5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_5; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2147 = 10'h6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_6; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2148 = 10'h7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_7; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2149 = 10'h8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_8; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2150 = 10'h9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_9; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2151 = 10'ha == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_10; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2152 = 10'hb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_11; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2153 = 10'hc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_12; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2154 = 10'hd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_13; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2155 = 10'he == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_14; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2156 = 10'hf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_15; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2157 = 10'h10 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_16; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2158 = 10'h11 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_17; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2159 = 10'h12 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_18; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2160 = 10'h13 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_19; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2161 = 10'h14 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_20; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2162 = 10'h15 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_21; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2163 = 10'h16 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_22; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2164 = 10'h17 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_23; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2165 = 10'h18 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_24; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2166 = 10'h19 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_25; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2167 = 10'h1a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_26; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2168 = 10'h1b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_27; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2169 = 10'h1c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_28; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2170 = 10'h1d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_29; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2171 = 10'h1e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_30; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2172 = 10'h1f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_31; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2173 = 10'h20 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_32; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2174 = 10'h21 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_33; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2175 = 10'h22 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_34; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2176 = 10'h23 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_35; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2177 = 10'h24 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_36; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2178 = 10'h25 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_37; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2179 = 10'h26 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_38; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2180 = 10'h27 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_39; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2181 = 10'h28 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_40; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2182 = 10'h29 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_41; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2183 = 10'h2a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_42; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2184 = 10'h2b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_43; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2185 = 10'h2c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_44; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2186 = 10'h2d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_45; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2187 = 10'h2e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_46; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2188 = 10'h2f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_47; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2189 = 10'h30 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_48; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2190 = 10'h31 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_49; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2191 = 10'h32 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_50; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2192 = 10'h33 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_51; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2193 = 10'h34 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_52; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2194 = 10'h35 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_53; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2195 = 10'h36 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_54; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2196 = 10'h37 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_55; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2197 = 10'h38 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_56; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2198 = 10'h39 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_57; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2199 = 10'h3a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_58; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2200 = 10'h3b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_59; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2201 = 10'h3c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_60; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2202 = 10'h3d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_61; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2203 = 10'h3e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_62; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2204 = 10'h3f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_63; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2205 = 10'h40 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_64; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2206 = 10'h41 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_65; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2207 = 10'h42 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_66; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2208 = 10'h43 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_67; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2209 = 10'h44 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_68; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2210 = 10'h45 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_69; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2211 = 10'h46 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_70; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2212 = 10'h47 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_71; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2213 = 10'h48 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_72; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2214 = 10'h49 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_73; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2215 = 10'h4a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_74; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2216 = 10'h4b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_75; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2217 = 10'h4c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_76; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2218 = 10'h4d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_77; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2219 = 10'h4e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_78; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2220 = 10'h4f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_79; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2221 = 10'h50 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_80; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2222 = 10'h51 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_81; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2223 = 10'h52 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_82; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2224 = 10'h53 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_83; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2225 = 10'h54 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_84; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2226 = 10'h55 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_85; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2227 = 10'h56 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_86; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2228 = 10'h57 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_87; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2229 = 10'h58 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_88; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2230 = 10'h59 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_89; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2231 = 10'h5a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_90; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2232 = 10'h5b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_91; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2233 = 10'h5c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_92; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2234 = 10'h5d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_93; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2235 = 10'h5e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_94; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2236 = 10'h5f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_95; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2237 = 10'h60 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_96; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2238 = 10'h61 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_97; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2239 = 10'h62 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_98; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2240 = 10'h63 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_99; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2241 = 10'h64 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_100; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2242 = 10'h65 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_101; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2243 = 10'h66 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_102; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2244 = 10'h67 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_103; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2245 = 10'h68 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_104; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2246 = 10'h69 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_105; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2247 = 10'h6a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_106; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2248 = 10'h6b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_107; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2249 = 10'h6c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_108; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2250 = 10'h6d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_109; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2251 = 10'h6e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_110; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2252 = 10'h6f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_111; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2253 = 10'h70 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_112; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2254 = 10'h71 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_113; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2255 = 10'h72 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_114; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2256 = 10'h73 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_115; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2257 = 10'h74 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_116; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2258 = 10'h75 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_117; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2259 = 10'h76 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_118; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2260 = 10'h77 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_119; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2261 = 10'h78 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_120; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2262 = 10'h79 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_121; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2263 = 10'h7a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_122; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2264 = 10'h7b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_123; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2265 = 10'h7c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_124; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2266 = 10'h7d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_125; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2267 = 10'h7e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_126; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2268 = 10'h7f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_127; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2269 = 10'h80 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_128; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2270 = 10'h81 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_129; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2271 = 10'h82 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_130; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2272 = 10'h83 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_131; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2273 = 10'h84 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_132; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2274 = 10'h85 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_133; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2275 = 10'h86 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_134; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2276 = 10'h87 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_135; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2277 = 10'h88 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_136; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2278 = 10'h89 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_137; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2279 = 10'h8a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_138; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2280 = 10'h8b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_139; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2281 = 10'h8c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_140; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2282 = 10'h8d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_141; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2283 = 10'h8e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_142; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2284 = 10'h8f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_143; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2285 = 10'h90 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_144; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2286 = 10'h91 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_145; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2287 = 10'h92 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_146; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2288 = 10'h93 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_147; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2289 = 10'h94 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_148; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2290 = 10'h95 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_149; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2291 = 10'h96 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_150; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2292 = 10'h97 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_151; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2293 = 10'h98 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_152; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2294 = 10'h99 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_153; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2295 = 10'h9a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_154; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2296 = 10'h9b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_155; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2297 = 10'h9c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_156; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2298 = 10'h9d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_157; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2299 = 10'h9e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_158; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2300 = 10'h9f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_159; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2301 = 10'ha0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_160; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2302 = 10'ha1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_161; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2303 = 10'ha2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_162; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2304 = 10'ha3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_163; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2305 = 10'ha4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_164; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2306 = 10'ha5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_165; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2307 = 10'ha6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_166; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2308 = 10'ha7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_167; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2309 = 10'ha8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_168; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2310 = 10'ha9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_169; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2311 = 10'haa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_170; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2312 = 10'hab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_171; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2313 = 10'hac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_172; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2314 = 10'had == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_173; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2315 = 10'hae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_174; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2316 = 10'haf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_175; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2317 = 10'hb0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_176; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2318 = 10'hb1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_177; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2319 = 10'hb2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_178; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2320 = 10'hb3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_179; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2321 = 10'hb4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_180; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2322 = 10'hb5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_181; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2323 = 10'hb6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_182; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2324 = 10'hb7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_183; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2325 = 10'hb8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_184; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2326 = 10'hb9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_185; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2327 = 10'hba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_186; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2328 = 10'hbb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_187; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2329 = 10'hbc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_188; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2330 = 10'hbd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_189; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2331 = 10'hbe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_190; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2332 = 10'hbf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_191; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2333 = 10'hc0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_192; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2334 = 10'hc1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_193; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2335 = 10'hc2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_194; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2336 = 10'hc3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_195; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2337 = 10'hc4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_196; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2338 = 10'hc5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_197; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2339 = 10'hc6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_198; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2340 = 10'hc7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_199; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2341 = 10'hc8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_200; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2342 = 10'hc9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_201; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2343 = 10'hca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_202; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2344 = 10'hcb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_203; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2345 = 10'hcc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_204; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2346 = 10'hcd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_205; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2347 = 10'hce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_206; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2348 = 10'hcf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_207; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2349 = 10'hd0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_208; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2350 = 10'hd1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_209; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2351 = 10'hd2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_210; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2352 = 10'hd3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_211; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2353 = 10'hd4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_212; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2354 = 10'hd5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_213; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2355 = 10'hd6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_214; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2356 = 10'hd7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_215; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2357 = 10'hd8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_216; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2358 = 10'hd9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_217; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2359 = 10'hda == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_218; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2360 = 10'hdb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_219; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2361 = 10'hdc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_220; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2362 = 10'hdd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_221; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2363 = 10'hde == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_222; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2364 = 10'hdf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_223; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2365 = 10'he0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_224; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2366 = 10'he1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_225; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2367 = 10'he2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_226; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2368 = 10'he3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_227; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2369 = 10'he4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_228; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2370 = 10'he5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_229; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2371 = 10'he6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_230; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2372 = 10'he7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_231; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2373 = 10'he8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_232; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2374 = 10'he9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_233; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2375 = 10'hea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_234; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2376 = 10'heb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_235; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2377 = 10'hec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_236; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2378 = 10'hed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_237; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2379 = 10'hee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_238; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2380 = 10'hef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_239; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2381 = 10'hf0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_240; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2382 = 10'hf1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_241; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2383 = 10'hf2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_242; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2384 = 10'hf3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_243; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2385 = 10'hf4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_244; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2386 = 10'hf5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_245; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2387 = 10'hf6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_246; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2388 = 10'hf7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_247; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2389 = 10'hf8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_248; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2390 = 10'hf9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_249; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2391 = 10'hfa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_250; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2392 = 10'hfb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_251; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2393 = 10'hfc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_252; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2394 = 10'hfd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_253; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2395 = 10'hfe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_254; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2396 = 10'hff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_255; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2397 = 10'h100 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_256; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2398 = 10'h101 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_257; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2399 = 10'h102 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_258; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2400 = 10'h103 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_259; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2401 = 10'h104 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_260; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2402 = 10'h105 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_261; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2403 = 10'h106 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_262; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2404 = 10'h107 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_263; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2405 = 10'h108 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_264; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2406 = 10'h109 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_265; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2407 = 10'h10a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_266; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2408 = 10'h10b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_267; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2409 = 10'h10c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_268; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2410 = 10'h10d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_269; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2411 = 10'h10e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_270; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2412 = 10'h10f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_271; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2413 = 10'h110 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_272; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2414 = 10'h111 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_273; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2415 = 10'h112 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_274; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2416 = 10'h113 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_275; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2417 = 10'h114 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_276; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2418 = 10'h115 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_277; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2419 = 10'h116 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_278; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2420 = 10'h117 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_279; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2421 = 10'h118 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_280; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2422 = 10'h119 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_281; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2423 = 10'h11a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_282; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2424 = 10'h11b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_283; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2425 = 10'h11c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_284; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2426 = 10'h11d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_285; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2427 = 10'h11e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_286; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2428 = 10'h11f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_287; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2429 = 10'h120 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_288; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2430 = 10'h121 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_289; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2431 = 10'h122 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_290; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2432 = 10'h123 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_291; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2433 = 10'h124 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_292; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2434 = 10'h125 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_293; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2435 = 10'h126 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_294; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2436 = 10'h127 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_295; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2437 = 10'h128 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_296; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2438 = 10'h129 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_297; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2439 = 10'h12a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_298; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2440 = 10'h12b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_299; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2441 = 10'h12c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_300; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2442 = 10'h12d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_301; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2443 = 10'h12e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_302; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2444 = 10'h12f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_303; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2445 = 10'h130 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_304; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2446 = 10'h131 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_305; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2447 = 10'h132 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_306; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2448 = 10'h133 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_307; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2449 = 10'h134 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_308; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2450 = 10'h135 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_309; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2451 = 10'h136 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_310; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2452 = 10'h137 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_311; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2453 = 10'h138 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_312; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2454 = 10'h139 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_313; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2455 = 10'h13a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_314; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2456 = 10'h13b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_315; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2457 = 10'h13c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_316; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2458 = 10'h13d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_317; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2459 = 10'h13e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_318; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2460 = 10'h13f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_319; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2461 = 10'h140 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_320; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2462 = 10'h141 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_321; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2463 = 10'h142 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_322; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2464 = 10'h143 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_323; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2465 = 10'h144 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_324; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2466 = 10'h145 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_325; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2467 = 10'h146 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_326; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2468 = 10'h147 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_327; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2469 = 10'h148 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_328; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2470 = 10'h149 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_329; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2471 = 10'h14a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_330; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2472 = 10'h14b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_331; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2473 = 10'h14c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_332; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2474 = 10'h14d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_333; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2475 = 10'h14e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_334; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2476 = 10'h14f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_335; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2477 = 10'h150 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_336; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2478 = 10'h151 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_337; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2479 = 10'h152 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_338; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2480 = 10'h153 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_339; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2481 = 10'h154 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_340; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2482 = 10'h155 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_341; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2483 = 10'h156 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_342; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2484 = 10'h157 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_343; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2485 = 10'h158 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_344; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2486 = 10'h159 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_345; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2487 = 10'h15a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_346; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2488 = 10'h15b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_347; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2489 = 10'h15c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_348; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2490 = 10'h15d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_349; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2491 = 10'h15e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_350; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2492 = 10'h15f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_351; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2493 = 10'h160 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_352; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2494 = 10'h161 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_353; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2495 = 10'h162 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_354; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2496 = 10'h163 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_355; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2497 = 10'h164 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_356; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2498 = 10'h165 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_357; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2499 = 10'h166 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_358; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2500 = 10'h167 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_359; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2501 = 10'h168 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_360; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2502 = 10'h169 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_361; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2503 = 10'h16a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_362; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2504 = 10'h16b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_363; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2505 = 10'h16c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_364; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2506 = 10'h16d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_365; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2507 = 10'h16e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_366; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2508 = 10'h16f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_367; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2509 = 10'h170 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_368; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2510 = 10'h171 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_369; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2511 = 10'h172 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_370; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2512 = 10'h173 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_371; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2513 = 10'h174 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_372; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2514 = 10'h175 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_373; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2515 = 10'h176 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_374; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2516 = 10'h177 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_375; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2517 = 10'h178 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_376; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2518 = 10'h179 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_377; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2519 = 10'h17a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_378; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2520 = 10'h17b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_379; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2521 = 10'h17c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_380; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2522 = 10'h17d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_381; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2523 = 10'h17e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_382; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2524 = 10'h17f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_383; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2525 = 10'h180 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_384; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2526 = 10'h181 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_385; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2527 = 10'h182 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_386; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2528 = 10'h183 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_387; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2529 = 10'h184 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_388; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2530 = 10'h185 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_389; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2531 = 10'h186 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_390; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2532 = 10'h187 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_391; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2533 = 10'h188 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_392; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2534 = 10'h189 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_393; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2535 = 10'h18a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_394; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2536 = 10'h18b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_395; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2537 = 10'h18c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_396; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2538 = 10'h18d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_397; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2539 = 10'h18e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_398; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2540 = 10'h18f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_399; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2541 = 10'h190 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_400; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2542 = 10'h191 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_401; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2543 = 10'h192 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_402; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2544 = 10'h193 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_403; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2545 = 10'h194 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_404; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2546 = 10'h195 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_405; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2547 = 10'h196 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_406; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2548 = 10'h197 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_407; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2549 = 10'h198 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_408; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2550 = 10'h199 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_409; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2551 = 10'h19a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_410; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2552 = 10'h19b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_411; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2553 = 10'h19c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_412; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2554 = 10'h19d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_413; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2555 = 10'h19e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_414; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2556 = 10'h19f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_415; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2557 = 10'h1a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_416; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2558 = 10'h1a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_417; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2559 = 10'h1a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_418; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2560 = 10'h1a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_419; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2561 = 10'h1a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_420; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2562 = 10'h1a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_421; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2563 = 10'h1a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_422; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2564 = 10'h1a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_423; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2565 = 10'h1a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_424; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2566 = 10'h1a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_425; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2567 = 10'h1aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_426; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2568 = 10'h1ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_427; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2569 = 10'h1ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_428; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2570 = 10'h1ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_429; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2571 = 10'h1ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_430; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2572 = 10'h1af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_431; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2573 = 10'h1b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_432; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2574 = 10'h1b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_433; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2575 = 10'h1b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_434; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2576 = 10'h1b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_435; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2577 = 10'h1b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_436; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2578 = 10'h1b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_437; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2579 = 10'h1b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_438; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2580 = 10'h1b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_439; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2581 = 10'h1b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_440; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2582 = 10'h1b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_441; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2583 = 10'h1ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_442; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2584 = 10'h1bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_443; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2585 = 10'h1bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_444; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2586 = 10'h1bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_445; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2587 = 10'h1be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_446; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2588 = 10'h1bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_447; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2589 = 10'h1c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_448; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2590 = 10'h1c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_449; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2591 = 10'h1c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_450; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2592 = 10'h1c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_451; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2593 = 10'h1c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_452; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2594 = 10'h1c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_453; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2595 = 10'h1c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_454; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2596 = 10'h1c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_455; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2597 = 10'h1c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_456; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2598 = 10'h1c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_457; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2599 = 10'h1ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_458; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2600 = 10'h1cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_459; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2601 = 10'h1cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_460; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2602 = 10'h1cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_461; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2603 = 10'h1ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_462; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2604 = 10'h1cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_463; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2605 = 10'h1d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_464; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2606 = 10'h1d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_465; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2607 = 10'h1d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_466; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2608 = 10'h1d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_467; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2609 = 10'h1d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_468; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2610 = 10'h1d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_469; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2611 = 10'h1d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_470; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2612 = 10'h1d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_471; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2613 = 10'h1d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_472; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2614 = 10'h1d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_473; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2615 = 10'h1da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_474; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2616 = 10'h1db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_475; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2617 = 10'h1dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_476; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2618 = 10'h1dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_477; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2619 = 10'h1de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_478; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2620 = 10'h1df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_479; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2621 = 10'h1e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_480; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2622 = 10'h1e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_481; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2623 = 10'h1e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_482; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2624 = 10'h1e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_483; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2625 = 10'h1e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_484; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2626 = 10'h1e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_485; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2627 = 10'h1e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_486; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2628 = 10'h1e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_487; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2629 = 10'h1e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_488; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2630 = 10'h1e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_489; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2631 = 10'h1ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_490; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2632 = 10'h1eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_491; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2633 = 10'h1ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_492; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2634 = 10'h1ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_493; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2635 = 10'h1ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_494; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2636 = 10'h1ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_495; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2637 = 10'h1f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_496; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2638 = 10'h1f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_497; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2639 = 10'h1f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_498; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2640 = 10'h1f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_499; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2641 = 10'h1f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_500; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2642 = 10'h1f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_501; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2643 = 10'h1f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_502; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2644 = 10'h1f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_503; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2645 = 10'h1f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_504; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2646 = 10'h1f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_505; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2647 = 10'h1fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_506; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2648 = 10'h1fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_507; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2649 = 10'h1fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_508; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2650 = 10'h1fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_509; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2651 = 10'h1fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_510; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2652 = 10'h1ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_511; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2653 = 10'h200 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_512; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2654 = 10'h201 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_513; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2655 = 10'h202 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_514; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2656 = 10'h203 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_515; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2657 = 10'h204 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_516; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2658 = 10'h205 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_517; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2659 = 10'h206 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_518; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2660 = 10'h207 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_519; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2661 = 10'h208 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_520; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2662 = 10'h209 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_521; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2663 = 10'h20a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_522; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2664 = 10'h20b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_523; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2665 = 10'h20c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_524; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2666 = 10'h20d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_525; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2667 = 10'h20e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_526; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2668 = 10'h20f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_527; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2669 = 10'h210 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_528; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2670 = 10'h211 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_529; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2671 = 10'h212 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_530; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2672 = 10'h213 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_531; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2673 = 10'h214 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_532; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2674 = 10'h215 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_533; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2675 = 10'h216 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_534; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2676 = 10'h217 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_535; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2677 = 10'h218 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_536; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2678 = 10'h219 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_537; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2679 = 10'h21a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_538; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2680 = 10'h21b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_539; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2681 = 10'h21c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_540; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2682 = 10'h21d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_541; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2683 = 10'h21e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_542; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2684 = 10'h21f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_543; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2685 = 10'h220 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_544; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2686 = 10'h221 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_545; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2687 = 10'h222 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_546; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2688 = 10'h223 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_547; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2689 = 10'h224 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_548; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2690 = 10'h225 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_549; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2691 = 10'h226 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_550; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2692 = 10'h227 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_551; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2693 = 10'h228 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_552; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2694 = 10'h229 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_553; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2695 = 10'h22a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_554; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2696 = 10'h22b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_555; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2697 = 10'h22c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_556; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2698 = 10'h22d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_557; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2699 = 10'h22e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_558; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2700 = 10'h22f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_559; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2701 = 10'h230 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_560; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2702 = 10'h231 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_561; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2703 = 10'h232 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_562; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2704 = 10'h233 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_563; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2705 = 10'h234 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_564; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2706 = 10'h235 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_565; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2707 = 10'h236 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_566; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2708 = 10'h237 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_567; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2709 = 10'h238 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_568; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2710 = 10'h239 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_569; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2711 = 10'h23a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_570; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2712 = 10'h23b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_571; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2713 = 10'h23c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_572; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2714 = 10'h23d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_573; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2715 = 10'h23e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_574; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2716 = 10'h23f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_575; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2717 = 10'h240 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_576; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2718 = 10'h241 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_577; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2719 = 10'h242 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_578; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2720 = 10'h243 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_579; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2721 = 10'h244 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_580; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2722 = 10'h245 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_581; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2723 = 10'h246 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_582; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2724 = 10'h247 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_583; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2725 = 10'h248 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_584; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2726 = 10'h249 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_585; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2727 = 10'h24a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_586; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2728 = 10'h24b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_587; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2729 = 10'h24c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_588; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2730 = 10'h24d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_589; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2731 = 10'h24e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_590; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2732 = 10'h24f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_591; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2733 = 10'h250 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_592; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2734 = 10'h251 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_593; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2735 = 10'h252 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_594; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2736 = 10'h253 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_595; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2737 = 10'h254 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_596; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2738 = 10'h255 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_597; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2739 = 10'h256 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_598; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2740 = 10'h257 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_599; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2741 = 10'h258 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_600; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2742 = 10'h259 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_601; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2743 = 10'h25a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_602; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2744 = 10'h25b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_603; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2745 = 10'h25c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_604; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2746 = 10'h25d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_605; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2747 = 10'h25e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_606; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2748 = 10'h25f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_607; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2749 = 10'h260 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_608; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2750 = 10'h261 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_609; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2751 = 10'h262 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_610; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2752 = 10'h263 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_611; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2753 = 10'h264 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_612; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2754 = 10'h265 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_613; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2755 = 10'h266 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_614; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2756 = 10'h267 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_615; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2757 = 10'h268 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_616; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2758 = 10'h269 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_617; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2759 = 10'h26a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_618; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2760 = 10'h26b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_619; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2761 = 10'h26c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_620; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2762 = 10'h26d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_621; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2763 = 10'h26e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_622; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2764 = 10'h26f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_623; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2765 = 10'h270 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_624; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2766 = 10'h271 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_625; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2767 = 10'h272 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_626; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2768 = 10'h273 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_627; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2769 = 10'h274 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_628; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2770 = 10'h275 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_629; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2771 = 10'h276 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_630; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2772 = 10'h277 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_631; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2773 = 10'h278 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_632; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2774 = 10'h279 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_633; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2775 = 10'h27a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_634; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2776 = 10'h27b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_635; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2777 = 10'h27c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_636; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2778 = 10'h27d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_637; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2779 = 10'h27e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_638; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2780 = 10'h27f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_639; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2781 = 10'h280 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_640; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2782 = 10'h281 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_641; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2783 = 10'h282 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_642; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2784 = 10'h283 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_643; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2785 = 10'h284 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_644; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2786 = 10'h285 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_645; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2787 = 10'h286 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_646; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2788 = 10'h287 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_647; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2789 = 10'h288 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_648; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2790 = 10'h289 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_649; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2791 = 10'h28a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_650; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2792 = 10'h28b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_651; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2793 = 10'h28c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_652; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2794 = 10'h28d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_653; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2795 = 10'h28e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_654; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2796 = 10'h28f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_655; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2797 = 10'h290 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_656; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2798 = 10'h291 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_657; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2799 = 10'h292 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_658; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2800 = 10'h293 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_659; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2801 = 10'h294 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_660; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2802 = 10'h295 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_661; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2803 = 10'h296 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_662; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2804 = 10'h297 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_663; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2805 = 10'h298 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_664; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2806 = 10'h299 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_665; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2807 = 10'h29a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_666; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2808 = 10'h29b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_667; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2809 = 10'h29c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_668; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2810 = 10'h29d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_669; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2811 = 10'h29e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_670; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2812 = 10'h29f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_671; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2813 = 10'h2a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_672; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2814 = 10'h2a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_673; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2815 = 10'h2a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_674; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2816 = 10'h2a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_675; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2817 = 10'h2a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_676; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2818 = 10'h2a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_677; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2819 = 10'h2a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_678; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2820 = 10'h2a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_679; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2821 = 10'h2a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_680; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2822 = 10'h2a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_681; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2823 = 10'h2aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_682; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2824 = 10'h2ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_683; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2825 = 10'h2ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_684; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2826 = 10'h2ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_685; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2827 = 10'h2ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_686; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2828 = 10'h2af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_687; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2829 = 10'h2b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_688; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2830 = 10'h2b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_689; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2831 = 10'h2b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_690; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2832 = 10'h2b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_691; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2833 = 10'h2b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_692; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2834 = 10'h2b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_693; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2835 = 10'h2b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_694; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2836 = 10'h2b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_695; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2837 = 10'h2b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_696; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2838 = 10'h2b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_697; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2839 = 10'h2ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_698; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2840 = 10'h2bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_699; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2841 = 10'h2bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_700; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2842 = 10'h2bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_701; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2843 = 10'h2be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_702; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2844 = 10'h2bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_703; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2845 = 10'h2c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_704; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2846 = 10'h2c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_705; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2847 = 10'h2c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_706; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2848 = 10'h2c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_707; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2849 = 10'h2c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_708; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2850 = 10'h2c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_709; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2851 = 10'h2c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_710; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2852 = 10'h2c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_711; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2853 = 10'h2c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_712; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2854 = 10'h2c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_713; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2855 = 10'h2ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_714; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2856 = 10'h2cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_715; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2857 = 10'h2cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_716; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2858 = 10'h2cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_717; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2859 = 10'h2ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_718; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2860 = 10'h2cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_719; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2861 = 10'h2d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_720; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2862 = 10'h2d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_721; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2863 = 10'h2d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_722; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2864 = 10'h2d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_723; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2865 = 10'h2d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_724; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2866 = 10'h2d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_725; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2867 = 10'h2d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_726; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2868 = 10'h2d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_727; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2869 = 10'h2d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_728; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2870 = 10'h2d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_729; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2871 = 10'h2da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_730; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2872 = 10'h2db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_731; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2873 = 10'h2dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_732; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2874 = 10'h2dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_733; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2875 = 10'h2de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_734; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2876 = 10'h2df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_735; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2877 = 10'h2e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_736; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2878 = 10'h2e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_737; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2879 = 10'h2e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_738; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2880 = 10'h2e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_739; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2881 = 10'h2e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_740; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2882 = 10'h2e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_741; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2883 = 10'h2e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_742; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2884 = 10'h2e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_743; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2885 = 10'h2e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_744; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2886 = 10'h2e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_745; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2887 = 10'h2ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_746; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2888 = 10'h2eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_747; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2889 = 10'h2ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_748; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2890 = 10'h2ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_749; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2891 = 10'h2ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_750; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2892 = 10'h2ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_751; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2893 = 10'h2f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_752; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2894 = 10'h2f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_753; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2895 = 10'h2f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_754; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2896 = 10'h2f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_755; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2897 = 10'h2f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_756; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2898 = 10'h2f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_757; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2899 = 10'h2f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_758; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2900 = 10'h2f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_759; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2901 = 10'h2f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_760; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2902 = 10'h2f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_761; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2903 = 10'h2fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_762; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2904 = 10'h2fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_763; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2905 = 10'h2fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_764; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2906 = 10'h2fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_765; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2907 = 10'h2fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_766; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2908 = 10'h2ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_767; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2909 = 10'h300 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_768; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2910 = 10'h301 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_769; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2911 = 10'h302 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_770; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2912 = 10'h303 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_771; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2913 = 10'h304 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_772; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2914 = 10'h305 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_773; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2915 = 10'h306 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_774; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2916 = 10'h307 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_775; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2917 = 10'h308 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_776; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2918 = 10'h309 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_777; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2919 = 10'h30a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_778; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2920 = 10'h30b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_779; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2921 = 10'h30c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_780; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2922 = 10'h30d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_781; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2923 = 10'h30e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_782; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2924 = 10'h30f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_783; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2925 = 10'h310 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_784; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2926 = 10'h311 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_785; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2927 = 10'h312 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_786; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2928 = 10'h313 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_787; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2929 = 10'h314 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_788; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2930 = 10'h315 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_789; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2931 = 10'h316 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_790; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2932 = 10'h317 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_791; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2933 = 10'h318 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_792; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2934 = 10'h319 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_793; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2935 = 10'h31a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_794; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2936 = 10'h31b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_795; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2937 = 10'h31c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_796; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2938 = 10'h31d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_797; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2939 = 10'h31e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_798; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2940 = 10'h31f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_799; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2941 = 10'h320 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_800; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2942 = 10'h321 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_801; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2943 = 10'h322 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_802; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2944 = 10'h323 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_803; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2945 = 10'h324 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_804; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2946 = 10'h325 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_805; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2947 = 10'h326 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_806; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2948 = 10'h327 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_807; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2949 = 10'h328 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_808; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2950 = 10'h329 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_809; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2951 = 10'h32a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_810; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2952 = 10'h32b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_811; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2953 = 10'h32c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_812; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2954 = 10'h32d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_813; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2955 = 10'h32e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_814; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2956 = 10'h32f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_815; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2957 = 10'h330 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_816; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2958 = 10'h331 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_817; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2959 = 10'h332 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_818; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2960 = 10'h333 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_819; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2961 = 10'h334 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_820; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2962 = 10'h335 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_821; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2963 = 10'h336 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_822; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2964 = 10'h337 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_823; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2965 = 10'h338 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_824; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2966 = 10'h339 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_825; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2967 = 10'h33a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_826; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2968 = 10'h33b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_827; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2969 = 10'h33c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_828; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2970 = 10'h33d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_829; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2971 = 10'h33e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_830; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2972 = 10'h33f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_831; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2973 = 10'h340 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_832; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2974 = 10'h341 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_833; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2975 = 10'h342 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_834; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2976 = 10'h343 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_835; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2977 = 10'h344 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_836; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2978 = 10'h345 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_837; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2979 = 10'h346 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_838; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2980 = 10'h347 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_839; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2981 = 10'h348 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_840; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2982 = 10'h349 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_841; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2983 = 10'h34a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_842; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2984 = 10'h34b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_843; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2985 = 10'h34c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_844; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2986 = 10'h34d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_845; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2987 = 10'h34e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_846; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2988 = 10'h34f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_847; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2989 = 10'h350 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_848; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2990 = 10'h351 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_849; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2991 = 10'h352 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_850; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2992 = 10'h353 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_851; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2993 = 10'h354 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_852; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2994 = 10'h355 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_853; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2995 = 10'h356 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_854; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2996 = 10'h357 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_855; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2997 = 10'h358 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_856; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2998 = 10'h359 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_857; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_2999 = 10'h35a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_858; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3000 = 10'h35b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_859; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3001 = 10'h35c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_860; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3002 = 10'h35d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_861; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3003 = 10'h35e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_862; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3004 = 10'h35f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_863; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3005 = 10'h360 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_864; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3006 = 10'h361 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_865; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3007 = 10'h362 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_866; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3008 = 10'h363 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_867; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3009 = 10'h364 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_868; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3010 = 10'h365 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_869; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3011 = 10'h366 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_870; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3012 = 10'h367 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_871; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3013 = 10'h368 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_872; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3014 = 10'h369 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_873; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3015 = 10'h36a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_874; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3016 = 10'h36b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_875; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3017 = 10'h36c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_876; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3018 = 10'h36d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_877; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3019 = 10'h36e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_878; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3020 = 10'h36f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_879; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3021 = 10'h370 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_880; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3022 = 10'h371 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_881; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3023 = 10'h372 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_882; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3024 = 10'h373 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_883; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3025 = 10'h374 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_884; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3026 = 10'h375 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_885; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3027 = 10'h376 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_886; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3028 = 10'h377 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_887; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3029 = 10'h378 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_888; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3030 = 10'h379 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_889; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3031 = 10'h37a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_890; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3032 = 10'h37b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_891; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3033 = 10'h37c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_892; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3034 = 10'h37d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_893; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3035 = 10'h37e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_894; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3036 = 10'h37f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_895; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3037 = 10'h380 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_896; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3038 = 10'h381 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_897; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3039 = 10'h382 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_898; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3040 = 10'h383 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_899; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3041 = 10'h384 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_900; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3042 = 10'h385 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_901; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3043 = 10'h386 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_902; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3044 = 10'h387 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_903; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3045 = 10'h388 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_904; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3046 = 10'h389 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_905; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3047 = 10'h38a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_906; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3048 = 10'h38b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_907; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3049 = 10'h38c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_908; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3050 = 10'h38d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_909; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3051 = 10'h38e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_910; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3052 = 10'h38f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_911; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3053 = 10'h390 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_912; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3054 = 10'h391 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_913; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3055 = 10'h392 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_914; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3056 = 10'h393 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_915; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3057 = 10'h394 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_916; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3058 = 10'h395 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_917; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3059 = 10'h396 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_918; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3060 = 10'h397 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_919; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3061 = 10'h398 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_920; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3062 = 10'h399 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_921; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3063 = 10'h39a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_922; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3064 = 10'h39b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_923; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3065 = 10'h39c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_924; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3066 = 10'h39d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_925; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3067 = 10'h39e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_926; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3068 = 10'h39f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_927; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3069 = 10'h3a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_928; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3070 = 10'h3a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_929; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3071 = 10'h3a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_930; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3072 = 10'h3a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_931; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3073 = 10'h3a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_932; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3074 = 10'h3a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_933; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3075 = 10'h3a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_934; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3076 = 10'h3a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_935; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3077 = 10'h3a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_936; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3078 = 10'h3a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_937; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3079 = 10'h3aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_938; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3080 = 10'h3ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_939; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3081 = 10'h3ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_940; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3082 = 10'h3ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_941; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3083 = 10'h3ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_942; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3084 = 10'h3af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_943; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3085 = 10'h3b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_944; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3086 = 10'h3b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_945; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3087 = 10'h3b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_946; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3088 = 10'h3b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_947; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3089 = 10'h3b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_948; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3090 = 10'h3b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_949; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3091 = 10'h3b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_950; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3092 = 10'h3b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_951; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3093 = 10'h3b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_952; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3094 = 10'h3b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_953; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3095 = 10'h3ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_954; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3096 = 10'h3bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_955; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3097 = 10'h3bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_956; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3098 = 10'h3bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_957; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3099 = 10'h3be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_958; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3100 = 10'h3bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_959; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3101 = 10'h3c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_960; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3102 = 10'h3c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_961; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3103 = 10'h3c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_962; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3104 = 10'h3c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_963; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3105 = 10'h3c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_964; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3106 = 10'h3c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_965; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3107 = 10'h3c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_966; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3108 = 10'h3c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_967; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3109 = 10'h3c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_968; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3110 = 10'h3c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_969; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3111 = 10'h3ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_970; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3112 = 10'h3cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_971; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3113 = 10'h3cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_972; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3114 = 10'h3cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_973; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3115 = 10'h3ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_974; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3116 = 10'h3cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_975; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3117 = 10'h3d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_976; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3118 = 10'h3d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_977; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3119 = 10'h3d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_978; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3120 = 10'h3d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_979; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3121 = 10'h3d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_980; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3122 = 10'h3d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_981; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3123 = 10'h3d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_982; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3124 = 10'h3d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_983; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3125 = 10'h3d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_984; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3126 = 10'h3d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_985; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3127 = 10'h3da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_986; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3128 = 10'h3db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_987; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3129 = 10'h3dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_988; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3130 = 10'h3dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_989; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3131 = 10'h3de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_990; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3132 = 10'h3df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_991; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3133 = 10'h3e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_992; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3134 = 10'h3e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_993; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3135 = 10'h3e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_994; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3136 = 10'h3e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_995; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3137 = 10'h3e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_996; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3138 = 10'h3e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_997; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3139 = 10'h3e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_998; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3140 = 10'h3e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_999; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3141 = 10'h3e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1000; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3142 = 10'h3e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1001; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3143 = 10'h3ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1002; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3144 = 10'h3eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1003; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3145 = 10'h3ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1004; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3146 = 10'h3ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1005; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3147 = 10'h3ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1006; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3148 = 10'h3ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1007; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3149 = 10'h3f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1008; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3150 = 10'h3f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1009; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3151 = 10'h3f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1010; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3152 = 10'h3f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1011; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3153 = 10'h3f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1012; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3154 = 10'h3f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1013; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3155 = 10'h3f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1014; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3156 = 10'h3f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1015; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3157 = 10'h3f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1016; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3158 = 10'h3f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1017; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3159 = 10'h3fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1018; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3160 = 10'h3fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1019; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3161 = 10'h3fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1020; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3162 = 10'h3fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1021; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3163 = 10'h3fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1022; // @[cpu.scala 201:{37,37} 46:20]
  wire [31:0] _GEN_3164 = 10'h3ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1023; // @[cpu.scala 201:{37,37} 46:20]
  assign io_rvfi_valid = 1'h0; // @[cpu.scala 219:17]
  assign io_rvfi_insn = MEMWBIR; // @[cpu.scala 218:16]
  assign io_rvfi_pc_rdata = CurPC; // @[cpu.scala 222:20]
  assign io_rvfi_pc_wdata = PC; // @[cpu.scala 224:20]
  assign io_rvfi_rs1_addr = io_rvfi_rst ? IFIDIR[19:15] : IFIDIR[19:15]; // @[cpu.scala 55:21 57:13 77:13]
  assign io_rvfi_rs2_addr = io_rvfi_rst ? IFIDIR[24:20] : IFIDIR[24:20]; // @[cpu.scala 55:21 58:13 78:13]
  assign io_rvfi_rs1_rdata = IDEXA; // @[cpu.scala 230:21]
  assign io_rvfi_rs2_rdata = IDEXB; // @[cpu.scala 232:21]
  assign io_rvfi_rd_addr = io_rvfi_rst ? MEMWBIR[11:7] : MEMWBIR[11:7]; // @[cpu.scala 55:21 63:13 83:13]
  assign io_rvfi_rd_wdata = MEMWBValue; // @[cpu.scala 215:20]
  assign io_rvfi_mem_addr = EXMEMALUOut[31:0]; // @[cpu.scala 236:20]
  assign io_rvfi_mem_rdata = MEMWBValue; // @[cpu.scala 238:21]
  assign io_rvfi_mem_wdata = {{32'd0}, DMemory_1}; // @[cpu.scala 240:21]
  assign io_rvfi_regs_0 = Regs_0; // @[cpu.scala 217:16]
  assign io_rvfi_regs_1 = Regs_1; // @[cpu.scala 217:16]
  assign io_rvfi_regs_2 = Regs_2; // @[cpu.scala 217:16]
  assign io_rvfi_regs_3 = Regs_3; // @[cpu.scala 217:16]
  assign io_rvfi_regs_4 = Regs_4; // @[cpu.scala 217:16]
  assign io_rvfi_regs_5 = Regs_5; // @[cpu.scala 217:16]
  assign io_rvfi_regs_6 = Regs_6; // @[cpu.scala 217:16]
  assign io_rvfi_regs_7 = Regs_7; // @[cpu.scala 217:16]
  assign io_rvfi_regs_8 = Regs_8; // @[cpu.scala 217:16]
  assign io_rvfi_regs_9 = Regs_9; // @[cpu.scala 217:16]
  assign io_rvfi_regs_10 = Regs_10; // @[cpu.scala 217:16]
  assign io_rvfi_regs_11 = Regs_11; // @[cpu.scala 217:16]
  assign io_rvfi_regs_12 = Regs_12; // @[cpu.scala 217:16]
  assign io_rvfi_regs_13 = Regs_13; // @[cpu.scala 217:16]
  assign io_rvfi_regs_14 = Regs_14; // @[cpu.scala 217:16]
  assign io_rvfi_regs_15 = Regs_15; // @[cpu.scala 217:16]
  assign io_rvfi_regs_16 = Regs_16; // @[cpu.scala 217:16]
  assign io_rvfi_regs_17 = Regs_17; // @[cpu.scala 217:16]
  assign io_rvfi_regs_18 = Regs_18; // @[cpu.scala 217:16]
  assign io_rvfi_regs_19 = Regs_19; // @[cpu.scala 217:16]
  assign io_rvfi_regs_20 = Regs_20; // @[cpu.scala 217:16]
  assign io_rvfi_regs_21 = Regs_21; // @[cpu.scala 217:16]
  assign io_rvfi_regs_22 = Regs_22; // @[cpu.scala 217:16]
  assign io_rvfi_regs_23 = Regs_23; // @[cpu.scala 217:16]
  assign io_rvfi_regs_24 = Regs_24; // @[cpu.scala 217:16]
  assign io_rvfi_regs_25 = Regs_25; // @[cpu.scala 217:16]
  assign io_rvfi_regs_26 = Regs_26; // @[cpu.scala 217:16]
  assign io_rvfi_regs_27 = Regs_27; // @[cpu.scala 217:16]
  assign io_rvfi_regs_28 = Regs_28; // @[cpu.scala 217:16]
  assign io_rvfi_regs_29 = Regs_29; // @[cpu.scala 217:16]
  assign io_rvfi_regs_30 = Regs_30; // @[cpu.scala 217:16]
  assign io_rvfi_regs_31 = Regs_31; // @[cpu.scala 217:16]
  always @(posedge clock) begin
    if (reset) begin // @[cpu.scala 42:19]
      PC <= 64'h0; // @[cpu.scala 42:19]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      if (~stall) begin // @[cpu.scala 117:27]
        if (~takeBranch) begin // @[cpu.scala 118:34]
          PC <= _PC_T_1; // @[cpu.scala 122:12]
        end else begin
          PC <= branchTarget; // @[cpu.scala 138:12]
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_0 <= io_rvfi_reg_data_in_0; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h0 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_0 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_1 <= io_rvfi_reg_data_in_1; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h1 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_1 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_2 <= io_rvfi_reg_data_in_2; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h2 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_2 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_3 <= io_rvfi_reg_data_in_3; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h3 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_3 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_4 <= io_rvfi_reg_data_in_4; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h4 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_4 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_5 <= io_rvfi_reg_data_in_5; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h5 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_5 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_6 <= io_rvfi_reg_data_in_6; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h6 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_6 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_7 <= io_rvfi_reg_data_in_7; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h7 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_7 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_8 <= io_rvfi_reg_data_in_8; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h8 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_8 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_9 <= io_rvfi_reg_data_in_9; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h9 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_9 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_10 <= io_rvfi_reg_data_in_10; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'ha == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_10 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_11 <= io_rvfi_reg_data_in_11; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'hb == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_11 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_12 <= io_rvfi_reg_data_in_12; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'hc == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_12 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_13 <= io_rvfi_reg_data_in_13; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'hd == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_13 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_14 <= io_rvfi_reg_data_in_14; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'he == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_14 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_15 <= io_rvfi_reg_data_in_15; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'hf == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_15 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_16 <= io_rvfi_reg_data_in_16; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h10 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_16 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_17 <= io_rvfi_reg_data_in_17; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h11 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_17 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_18 <= io_rvfi_reg_data_in_18; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h12 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_18 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_19 <= io_rvfi_reg_data_in_19; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h13 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_19 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_20 <= io_rvfi_reg_data_in_20; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h14 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_20 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_21 <= io_rvfi_reg_data_in_21; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h15 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_21 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_22 <= io_rvfi_reg_data_in_22; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h16 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_22 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_23 <= io_rvfi_reg_data_in_23; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h17 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_23 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_24 <= io_rvfi_reg_data_in_24; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h18 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_24 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_25 <= io_rvfi_reg_data_in_25; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h19 == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_25 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_26 <= io_rvfi_reg_data_in_26; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h1a == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_26 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_27 <= io_rvfi_reg_data_in_27; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h1b == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_27 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_28 <= io_rvfi_reg_data_in_28; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h1c == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_28 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_29 <= io_rvfi_reg_data_in_29; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h1d == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_29 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_30 <= io_rvfi_reg_data_in_30; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h1e == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_30 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      Regs_31 <= io_rvfi_reg_data_in_31; // @[cpu.scala 68:14]
    end else if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 210:74]
      if (5'h1f == MEMWBrd) begin // @[cpu.scala 211:21]
        Regs_31 <= MEMWBValue; // @[cpu.scala 211:21]
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      if (~stall) begin // @[cpu.scala 117:27]
        if (bypassAFromEX) begin // @[cpu.scala 144:27]
          IDEXA <= _A_T_1; // @[cpu.scala 146:11]
        end else if (bypassAFromMEM) begin // @[cpu.scala 147:34]
          IDEXA <= EXMEMALUOut; // @[cpu.scala 149:11]
        end else begin
          IDEXA <= _GEN_1061;
        end
      end else begin
        IDEXA <= 64'h0;
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      if (~stall) begin // @[cpu.scala 117:27]
        if (bypassBFromEX) begin // @[cpu.scala 157:27]
          IDEXB <= _B_T_1; // @[cpu.scala 159:11]
        end else if (bypassBFromMEM) begin // @[cpu.scala 160:34]
          IDEXB <= EXMEMALUOut; // @[cpu.scala 162:11]
        end else begin
          IDEXB <= _GEN_1099;
        end
      end else begin
        IDEXB <= 64'h0;
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      EXMEMB <= IDEXB; // @[cpu.scala 193:12]
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      if (_stall_T_9) begin // @[cpu.scala 178:25]
        EXMEMALUOut <= _EXMEMALUOut_T_6; // @[cpu.scala 179:19]
      end else if (IDEXop == 7'h23) begin // @[cpu.scala 180:31]
        EXMEMALUOut <= _EXMEMALUOut_T_15; // @[cpu.scala 181:19]
      end else if (_bypassAFromEX_T_3) begin // @[cpu.scala 185:34]
        EXMEMALUOut <= _A_T_1; // @[cpu.scala 188:19]
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      if (_bypassAFromMEM_T_3) begin // @[cpu.scala 196:29]
        MEMWBValue <= EXMEMALUOut; // @[cpu.scala 197:18]
      end else if (_stall_T) begin // @[cpu.scala 198:32]
        MEMWBValue <= {{32'd0}, _GEN_2140}; // @[cpu.scala 199:18]
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_0 <= io_rvfi_mem_data_in_0; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_0 <= _GEN_2141;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1 <= io_rvfi_mem_data_in_1; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1 <= _GEN_2142;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_2 <= io_rvfi_mem_data_in_2; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_2 <= _GEN_2143;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_3 <= io_rvfi_mem_data_in_3; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_3 <= _GEN_2144;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_4 <= io_rvfi_mem_data_in_4; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_4 <= _GEN_2145;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_5 <= io_rvfi_mem_data_in_5; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_5 <= _GEN_2146;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_6 <= io_rvfi_mem_data_in_6; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_6 <= _GEN_2147;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_7 <= io_rvfi_mem_data_in_7; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_7 <= _GEN_2148;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_8 <= io_rvfi_mem_data_in_8; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_8 <= _GEN_2149;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_9 <= io_rvfi_mem_data_in_9; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_9 <= _GEN_2150;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_10 <= io_rvfi_mem_data_in_10; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_10 <= _GEN_2151;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_11 <= io_rvfi_mem_data_in_11; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_11 <= _GEN_2152;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_12 <= io_rvfi_mem_data_in_12; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_12 <= _GEN_2153;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_13 <= io_rvfi_mem_data_in_13; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_13 <= _GEN_2154;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_14 <= io_rvfi_mem_data_in_14; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_14 <= _GEN_2155;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_15 <= io_rvfi_mem_data_in_15; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_15 <= _GEN_2156;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_16 <= io_rvfi_mem_data_in_16; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_16 <= _GEN_2157;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_17 <= io_rvfi_mem_data_in_17; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_17 <= _GEN_2158;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_18 <= io_rvfi_mem_data_in_18; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_18 <= _GEN_2159;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_19 <= io_rvfi_mem_data_in_19; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_19 <= _GEN_2160;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_20 <= io_rvfi_mem_data_in_20; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_20 <= _GEN_2161;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_21 <= io_rvfi_mem_data_in_21; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_21 <= _GEN_2162;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_22 <= io_rvfi_mem_data_in_22; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_22 <= _GEN_2163;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_23 <= io_rvfi_mem_data_in_23; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_23 <= _GEN_2164;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_24 <= io_rvfi_mem_data_in_24; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_24 <= _GEN_2165;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_25 <= io_rvfi_mem_data_in_25; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_25 <= _GEN_2166;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_26 <= io_rvfi_mem_data_in_26; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_26 <= _GEN_2167;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_27 <= io_rvfi_mem_data_in_27; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_27 <= _GEN_2168;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_28 <= io_rvfi_mem_data_in_28; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_28 <= _GEN_2169;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_29 <= io_rvfi_mem_data_in_29; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_29 <= _GEN_2170;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_30 <= io_rvfi_mem_data_in_30; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_30 <= _GEN_2171;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_31 <= io_rvfi_mem_data_in_31; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_31 <= _GEN_2172;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_32 <= io_rvfi_mem_data_in_32; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_32 <= _GEN_2173;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_33 <= io_rvfi_mem_data_in_33; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_33 <= _GEN_2174;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_34 <= io_rvfi_mem_data_in_34; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_34 <= _GEN_2175;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_35 <= io_rvfi_mem_data_in_35; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_35 <= _GEN_2176;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_36 <= io_rvfi_mem_data_in_36; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_36 <= _GEN_2177;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_37 <= io_rvfi_mem_data_in_37; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_37 <= _GEN_2178;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_38 <= io_rvfi_mem_data_in_38; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_38 <= _GEN_2179;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_39 <= io_rvfi_mem_data_in_39; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_39 <= _GEN_2180;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_40 <= io_rvfi_mem_data_in_40; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_40 <= _GEN_2181;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_41 <= io_rvfi_mem_data_in_41; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_41 <= _GEN_2182;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_42 <= io_rvfi_mem_data_in_42; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_42 <= _GEN_2183;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_43 <= io_rvfi_mem_data_in_43; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_43 <= _GEN_2184;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_44 <= io_rvfi_mem_data_in_44; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_44 <= _GEN_2185;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_45 <= io_rvfi_mem_data_in_45; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_45 <= _GEN_2186;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_46 <= io_rvfi_mem_data_in_46; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_46 <= _GEN_2187;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_47 <= io_rvfi_mem_data_in_47; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_47 <= _GEN_2188;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_48 <= io_rvfi_mem_data_in_48; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_48 <= _GEN_2189;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_49 <= io_rvfi_mem_data_in_49; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_49 <= _GEN_2190;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_50 <= io_rvfi_mem_data_in_50; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_50 <= _GEN_2191;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_51 <= io_rvfi_mem_data_in_51; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_51 <= _GEN_2192;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_52 <= io_rvfi_mem_data_in_52; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_52 <= _GEN_2193;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_53 <= io_rvfi_mem_data_in_53; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_53 <= _GEN_2194;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_54 <= io_rvfi_mem_data_in_54; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_54 <= _GEN_2195;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_55 <= io_rvfi_mem_data_in_55; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_55 <= _GEN_2196;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_56 <= io_rvfi_mem_data_in_56; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_56 <= _GEN_2197;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_57 <= io_rvfi_mem_data_in_57; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_57 <= _GEN_2198;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_58 <= io_rvfi_mem_data_in_58; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_58 <= _GEN_2199;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_59 <= io_rvfi_mem_data_in_59; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_59 <= _GEN_2200;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_60 <= io_rvfi_mem_data_in_60; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_60 <= _GEN_2201;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_61 <= io_rvfi_mem_data_in_61; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_61 <= _GEN_2202;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_62 <= io_rvfi_mem_data_in_62; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_62 <= _GEN_2203;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_63 <= io_rvfi_mem_data_in_63; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_63 <= _GEN_2204;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_64 <= io_rvfi_mem_data_in_64; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_64 <= _GEN_2205;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_65 <= io_rvfi_mem_data_in_65; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_65 <= _GEN_2206;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_66 <= io_rvfi_mem_data_in_66; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_66 <= _GEN_2207;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_67 <= io_rvfi_mem_data_in_67; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_67 <= _GEN_2208;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_68 <= io_rvfi_mem_data_in_68; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_68 <= _GEN_2209;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_69 <= io_rvfi_mem_data_in_69; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_69 <= _GEN_2210;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_70 <= io_rvfi_mem_data_in_70; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_70 <= _GEN_2211;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_71 <= io_rvfi_mem_data_in_71; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_71 <= _GEN_2212;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_72 <= io_rvfi_mem_data_in_72; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_72 <= _GEN_2213;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_73 <= io_rvfi_mem_data_in_73; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_73 <= _GEN_2214;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_74 <= io_rvfi_mem_data_in_74; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_74 <= _GEN_2215;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_75 <= io_rvfi_mem_data_in_75; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_75 <= _GEN_2216;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_76 <= io_rvfi_mem_data_in_76; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_76 <= _GEN_2217;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_77 <= io_rvfi_mem_data_in_77; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_77 <= _GEN_2218;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_78 <= io_rvfi_mem_data_in_78; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_78 <= _GEN_2219;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_79 <= io_rvfi_mem_data_in_79; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_79 <= _GEN_2220;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_80 <= io_rvfi_mem_data_in_80; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_80 <= _GEN_2221;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_81 <= io_rvfi_mem_data_in_81; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_81 <= _GEN_2222;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_82 <= io_rvfi_mem_data_in_82; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_82 <= _GEN_2223;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_83 <= io_rvfi_mem_data_in_83; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_83 <= _GEN_2224;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_84 <= io_rvfi_mem_data_in_84; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_84 <= _GEN_2225;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_85 <= io_rvfi_mem_data_in_85; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_85 <= _GEN_2226;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_86 <= io_rvfi_mem_data_in_86; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_86 <= _GEN_2227;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_87 <= io_rvfi_mem_data_in_87; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_87 <= _GEN_2228;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_88 <= io_rvfi_mem_data_in_88; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_88 <= _GEN_2229;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_89 <= io_rvfi_mem_data_in_89; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_89 <= _GEN_2230;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_90 <= io_rvfi_mem_data_in_90; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_90 <= _GEN_2231;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_91 <= io_rvfi_mem_data_in_91; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_91 <= _GEN_2232;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_92 <= io_rvfi_mem_data_in_92; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_92 <= _GEN_2233;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_93 <= io_rvfi_mem_data_in_93; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_93 <= _GEN_2234;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_94 <= io_rvfi_mem_data_in_94; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_94 <= _GEN_2235;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_95 <= io_rvfi_mem_data_in_95; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_95 <= _GEN_2236;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_96 <= io_rvfi_mem_data_in_96; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_96 <= _GEN_2237;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_97 <= io_rvfi_mem_data_in_97; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_97 <= _GEN_2238;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_98 <= io_rvfi_mem_data_in_98; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_98 <= _GEN_2239;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_99 <= io_rvfi_mem_data_in_99; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_99 <= _GEN_2240;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_100 <= io_rvfi_mem_data_in_100; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_100 <= _GEN_2241;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_101 <= io_rvfi_mem_data_in_101; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_101 <= _GEN_2242;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_102 <= io_rvfi_mem_data_in_102; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_102 <= _GEN_2243;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_103 <= io_rvfi_mem_data_in_103; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_103 <= _GEN_2244;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_104 <= io_rvfi_mem_data_in_104; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_104 <= _GEN_2245;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_105 <= io_rvfi_mem_data_in_105; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_105 <= _GEN_2246;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_106 <= io_rvfi_mem_data_in_106; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_106 <= _GEN_2247;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_107 <= io_rvfi_mem_data_in_107; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_107 <= _GEN_2248;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_108 <= io_rvfi_mem_data_in_108; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_108 <= _GEN_2249;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_109 <= io_rvfi_mem_data_in_109; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_109 <= _GEN_2250;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_110 <= io_rvfi_mem_data_in_110; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_110 <= _GEN_2251;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_111 <= io_rvfi_mem_data_in_111; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_111 <= _GEN_2252;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_112 <= io_rvfi_mem_data_in_112; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_112 <= _GEN_2253;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_113 <= io_rvfi_mem_data_in_113; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_113 <= _GEN_2254;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_114 <= io_rvfi_mem_data_in_114; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_114 <= _GEN_2255;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_115 <= io_rvfi_mem_data_in_115; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_115 <= _GEN_2256;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_116 <= io_rvfi_mem_data_in_116; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_116 <= _GEN_2257;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_117 <= io_rvfi_mem_data_in_117; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_117 <= _GEN_2258;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_118 <= io_rvfi_mem_data_in_118; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_118 <= _GEN_2259;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_119 <= io_rvfi_mem_data_in_119; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_119 <= _GEN_2260;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_120 <= io_rvfi_mem_data_in_120; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_120 <= _GEN_2261;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_121 <= io_rvfi_mem_data_in_121; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_121 <= _GEN_2262;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_122 <= io_rvfi_mem_data_in_122; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_122 <= _GEN_2263;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_123 <= io_rvfi_mem_data_in_123; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_123 <= _GEN_2264;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_124 <= io_rvfi_mem_data_in_124; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_124 <= _GEN_2265;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_125 <= io_rvfi_mem_data_in_125; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_125 <= _GEN_2266;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_126 <= io_rvfi_mem_data_in_126; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_126 <= _GEN_2267;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_127 <= io_rvfi_mem_data_in_127; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_127 <= _GEN_2268;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_128 <= io_rvfi_mem_data_in_128; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_128 <= _GEN_2269;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_129 <= io_rvfi_mem_data_in_129; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_129 <= _GEN_2270;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_130 <= io_rvfi_mem_data_in_130; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_130 <= _GEN_2271;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_131 <= io_rvfi_mem_data_in_131; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_131 <= _GEN_2272;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_132 <= io_rvfi_mem_data_in_132; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_132 <= _GEN_2273;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_133 <= io_rvfi_mem_data_in_133; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_133 <= _GEN_2274;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_134 <= io_rvfi_mem_data_in_134; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_134 <= _GEN_2275;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_135 <= io_rvfi_mem_data_in_135; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_135 <= _GEN_2276;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_136 <= io_rvfi_mem_data_in_136; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_136 <= _GEN_2277;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_137 <= io_rvfi_mem_data_in_137; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_137 <= _GEN_2278;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_138 <= io_rvfi_mem_data_in_138; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_138 <= _GEN_2279;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_139 <= io_rvfi_mem_data_in_139; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_139 <= _GEN_2280;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_140 <= io_rvfi_mem_data_in_140; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_140 <= _GEN_2281;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_141 <= io_rvfi_mem_data_in_141; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_141 <= _GEN_2282;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_142 <= io_rvfi_mem_data_in_142; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_142 <= _GEN_2283;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_143 <= io_rvfi_mem_data_in_143; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_143 <= _GEN_2284;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_144 <= io_rvfi_mem_data_in_144; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_144 <= _GEN_2285;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_145 <= io_rvfi_mem_data_in_145; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_145 <= _GEN_2286;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_146 <= io_rvfi_mem_data_in_146; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_146 <= _GEN_2287;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_147 <= io_rvfi_mem_data_in_147; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_147 <= _GEN_2288;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_148 <= io_rvfi_mem_data_in_148; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_148 <= _GEN_2289;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_149 <= io_rvfi_mem_data_in_149; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_149 <= _GEN_2290;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_150 <= io_rvfi_mem_data_in_150; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_150 <= _GEN_2291;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_151 <= io_rvfi_mem_data_in_151; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_151 <= _GEN_2292;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_152 <= io_rvfi_mem_data_in_152; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_152 <= _GEN_2293;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_153 <= io_rvfi_mem_data_in_153; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_153 <= _GEN_2294;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_154 <= io_rvfi_mem_data_in_154; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_154 <= _GEN_2295;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_155 <= io_rvfi_mem_data_in_155; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_155 <= _GEN_2296;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_156 <= io_rvfi_mem_data_in_156; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_156 <= _GEN_2297;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_157 <= io_rvfi_mem_data_in_157; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_157 <= _GEN_2298;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_158 <= io_rvfi_mem_data_in_158; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_158 <= _GEN_2299;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_159 <= io_rvfi_mem_data_in_159; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_159 <= _GEN_2300;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_160 <= io_rvfi_mem_data_in_160; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_160 <= _GEN_2301;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_161 <= io_rvfi_mem_data_in_161; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_161 <= _GEN_2302;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_162 <= io_rvfi_mem_data_in_162; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_162 <= _GEN_2303;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_163 <= io_rvfi_mem_data_in_163; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_163 <= _GEN_2304;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_164 <= io_rvfi_mem_data_in_164; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_164 <= _GEN_2305;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_165 <= io_rvfi_mem_data_in_165; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_165 <= _GEN_2306;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_166 <= io_rvfi_mem_data_in_166; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_166 <= _GEN_2307;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_167 <= io_rvfi_mem_data_in_167; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_167 <= _GEN_2308;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_168 <= io_rvfi_mem_data_in_168; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_168 <= _GEN_2309;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_169 <= io_rvfi_mem_data_in_169; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_169 <= _GEN_2310;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_170 <= io_rvfi_mem_data_in_170; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_170 <= _GEN_2311;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_171 <= io_rvfi_mem_data_in_171; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_171 <= _GEN_2312;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_172 <= io_rvfi_mem_data_in_172; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_172 <= _GEN_2313;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_173 <= io_rvfi_mem_data_in_173; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_173 <= _GEN_2314;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_174 <= io_rvfi_mem_data_in_174; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_174 <= _GEN_2315;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_175 <= io_rvfi_mem_data_in_175; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_175 <= _GEN_2316;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_176 <= io_rvfi_mem_data_in_176; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_176 <= _GEN_2317;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_177 <= io_rvfi_mem_data_in_177; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_177 <= _GEN_2318;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_178 <= io_rvfi_mem_data_in_178; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_178 <= _GEN_2319;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_179 <= io_rvfi_mem_data_in_179; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_179 <= _GEN_2320;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_180 <= io_rvfi_mem_data_in_180; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_180 <= _GEN_2321;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_181 <= io_rvfi_mem_data_in_181; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_181 <= _GEN_2322;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_182 <= io_rvfi_mem_data_in_182; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_182 <= _GEN_2323;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_183 <= io_rvfi_mem_data_in_183; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_183 <= _GEN_2324;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_184 <= io_rvfi_mem_data_in_184; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_184 <= _GEN_2325;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_185 <= io_rvfi_mem_data_in_185; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_185 <= _GEN_2326;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_186 <= io_rvfi_mem_data_in_186; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_186 <= _GEN_2327;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_187 <= io_rvfi_mem_data_in_187; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_187 <= _GEN_2328;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_188 <= io_rvfi_mem_data_in_188; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_188 <= _GEN_2329;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_189 <= io_rvfi_mem_data_in_189; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_189 <= _GEN_2330;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_190 <= io_rvfi_mem_data_in_190; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_190 <= _GEN_2331;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_191 <= io_rvfi_mem_data_in_191; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_191 <= _GEN_2332;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_192 <= io_rvfi_mem_data_in_192; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_192 <= _GEN_2333;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_193 <= io_rvfi_mem_data_in_193; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_193 <= _GEN_2334;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_194 <= io_rvfi_mem_data_in_194; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_194 <= _GEN_2335;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_195 <= io_rvfi_mem_data_in_195; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_195 <= _GEN_2336;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_196 <= io_rvfi_mem_data_in_196; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_196 <= _GEN_2337;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_197 <= io_rvfi_mem_data_in_197; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_197 <= _GEN_2338;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_198 <= io_rvfi_mem_data_in_198; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_198 <= _GEN_2339;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_199 <= io_rvfi_mem_data_in_199; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_199 <= _GEN_2340;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_200 <= io_rvfi_mem_data_in_200; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_200 <= _GEN_2341;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_201 <= io_rvfi_mem_data_in_201; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_201 <= _GEN_2342;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_202 <= io_rvfi_mem_data_in_202; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_202 <= _GEN_2343;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_203 <= io_rvfi_mem_data_in_203; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_203 <= _GEN_2344;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_204 <= io_rvfi_mem_data_in_204; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_204 <= _GEN_2345;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_205 <= io_rvfi_mem_data_in_205; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_205 <= _GEN_2346;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_206 <= io_rvfi_mem_data_in_206; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_206 <= _GEN_2347;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_207 <= io_rvfi_mem_data_in_207; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_207 <= _GEN_2348;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_208 <= io_rvfi_mem_data_in_208; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_208 <= _GEN_2349;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_209 <= io_rvfi_mem_data_in_209; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_209 <= _GEN_2350;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_210 <= io_rvfi_mem_data_in_210; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_210 <= _GEN_2351;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_211 <= io_rvfi_mem_data_in_211; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_211 <= _GEN_2352;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_212 <= io_rvfi_mem_data_in_212; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_212 <= _GEN_2353;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_213 <= io_rvfi_mem_data_in_213; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_213 <= _GEN_2354;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_214 <= io_rvfi_mem_data_in_214; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_214 <= _GEN_2355;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_215 <= io_rvfi_mem_data_in_215; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_215 <= _GEN_2356;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_216 <= io_rvfi_mem_data_in_216; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_216 <= _GEN_2357;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_217 <= io_rvfi_mem_data_in_217; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_217 <= _GEN_2358;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_218 <= io_rvfi_mem_data_in_218; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_218 <= _GEN_2359;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_219 <= io_rvfi_mem_data_in_219; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_219 <= _GEN_2360;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_220 <= io_rvfi_mem_data_in_220; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_220 <= _GEN_2361;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_221 <= io_rvfi_mem_data_in_221; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_221 <= _GEN_2362;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_222 <= io_rvfi_mem_data_in_222; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_222 <= _GEN_2363;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_223 <= io_rvfi_mem_data_in_223; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_223 <= _GEN_2364;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_224 <= io_rvfi_mem_data_in_224; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_224 <= _GEN_2365;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_225 <= io_rvfi_mem_data_in_225; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_225 <= _GEN_2366;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_226 <= io_rvfi_mem_data_in_226; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_226 <= _GEN_2367;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_227 <= io_rvfi_mem_data_in_227; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_227 <= _GEN_2368;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_228 <= io_rvfi_mem_data_in_228; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_228 <= _GEN_2369;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_229 <= io_rvfi_mem_data_in_229; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_229 <= _GEN_2370;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_230 <= io_rvfi_mem_data_in_230; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_230 <= _GEN_2371;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_231 <= io_rvfi_mem_data_in_231; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_231 <= _GEN_2372;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_232 <= io_rvfi_mem_data_in_232; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_232 <= _GEN_2373;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_233 <= io_rvfi_mem_data_in_233; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_233 <= _GEN_2374;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_234 <= io_rvfi_mem_data_in_234; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_234 <= _GEN_2375;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_235 <= io_rvfi_mem_data_in_235; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_235 <= _GEN_2376;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_236 <= io_rvfi_mem_data_in_236; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_236 <= _GEN_2377;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_237 <= io_rvfi_mem_data_in_237; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_237 <= _GEN_2378;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_238 <= io_rvfi_mem_data_in_238; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_238 <= _GEN_2379;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_239 <= io_rvfi_mem_data_in_239; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_239 <= _GEN_2380;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_240 <= io_rvfi_mem_data_in_240; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_240 <= _GEN_2381;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_241 <= io_rvfi_mem_data_in_241; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_241 <= _GEN_2382;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_242 <= io_rvfi_mem_data_in_242; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_242 <= _GEN_2383;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_243 <= io_rvfi_mem_data_in_243; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_243 <= _GEN_2384;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_244 <= io_rvfi_mem_data_in_244; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_244 <= _GEN_2385;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_245 <= io_rvfi_mem_data_in_245; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_245 <= _GEN_2386;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_246 <= io_rvfi_mem_data_in_246; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_246 <= _GEN_2387;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_247 <= io_rvfi_mem_data_in_247; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_247 <= _GEN_2388;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_248 <= io_rvfi_mem_data_in_248; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_248 <= _GEN_2389;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_249 <= io_rvfi_mem_data_in_249; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_249 <= _GEN_2390;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_250 <= io_rvfi_mem_data_in_250; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_250 <= _GEN_2391;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_251 <= io_rvfi_mem_data_in_251; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_251 <= _GEN_2392;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_252 <= io_rvfi_mem_data_in_252; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_252 <= _GEN_2393;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_253 <= io_rvfi_mem_data_in_253; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_253 <= _GEN_2394;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_254 <= io_rvfi_mem_data_in_254; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_254 <= _GEN_2395;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_255 <= io_rvfi_mem_data_in_255; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_255 <= _GEN_2396;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_256 <= io_rvfi_mem_data_in_256; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_256 <= _GEN_2397;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_257 <= io_rvfi_mem_data_in_257; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_257 <= _GEN_2398;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_258 <= io_rvfi_mem_data_in_258; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_258 <= _GEN_2399;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_259 <= io_rvfi_mem_data_in_259; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_259 <= _GEN_2400;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_260 <= io_rvfi_mem_data_in_260; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_260 <= _GEN_2401;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_261 <= io_rvfi_mem_data_in_261; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_261 <= _GEN_2402;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_262 <= io_rvfi_mem_data_in_262; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_262 <= _GEN_2403;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_263 <= io_rvfi_mem_data_in_263; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_263 <= _GEN_2404;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_264 <= io_rvfi_mem_data_in_264; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_264 <= _GEN_2405;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_265 <= io_rvfi_mem_data_in_265; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_265 <= _GEN_2406;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_266 <= io_rvfi_mem_data_in_266; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_266 <= _GEN_2407;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_267 <= io_rvfi_mem_data_in_267; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_267 <= _GEN_2408;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_268 <= io_rvfi_mem_data_in_268; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_268 <= _GEN_2409;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_269 <= io_rvfi_mem_data_in_269; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_269 <= _GEN_2410;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_270 <= io_rvfi_mem_data_in_270; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_270 <= _GEN_2411;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_271 <= io_rvfi_mem_data_in_271; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_271 <= _GEN_2412;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_272 <= io_rvfi_mem_data_in_272; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_272 <= _GEN_2413;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_273 <= io_rvfi_mem_data_in_273; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_273 <= _GEN_2414;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_274 <= io_rvfi_mem_data_in_274; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_274 <= _GEN_2415;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_275 <= io_rvfi_mem_data_in_275; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_275 <= _GEN_2416;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_276 <= io_rvfi_mem_data_in_276; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_276 <= _GEN_2417;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_277 <= io_rvfi_mem_data_in_277; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_277 <= _GEN_2418;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_278 <= io_rvfi_mem_data_in_278; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_278 <= _GEN_2419;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_279 <= io_rvfi_mem_data_in_279; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_279 <= _GEN_2420;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_280 <= io_rvfi_mem_data_in_280; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_280 <= _GEN_2421;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_281 <= io_rvfi_mem_data_in_281; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_281 <= _GEN_2422;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_282 <= io_rvfi_mem_data_in_282; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_282 <= _GEN_2423;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_283 <= io_rvfi_mem_data_in_283; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_283 <= _GEN_2424;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_284 <= io_rvfi_mem_data_in_284; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_284 <= _GEN_2425;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_285 <= io_rvfi_mem_data_in_285; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_285 <= _GEN_2426;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_286 <= io_rvfi_mem_data_in_286; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_286 <= _GEN_2427;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_287 <= io_rvfi_mem_data_in_287; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_287 <= _GEN_2428;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_288 <= io_rvfi_mem_data_in_288; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_288 <= _GEN_2429;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_289 <= io_rvfi_mem_data_in_289; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_289 <= _GEN_2430;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_290 <= io_rvfi_mem_data_in_290; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_290 <= _GEN_2431;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_291 <= io_rvfi_mem_data_in_291; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_291 <= _GEN_2432;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_292 <= io_rvfi_mem_data_in_292; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_292 <= _GEN_2433;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_293 <= io_rvfi_mem_data_in_293; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_293 <= _GEN_2434;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_294 <= io_rvfi_mem_data_in_294; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_294 <= _GEN_2435;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_295 <= io_rvfi_mem_data_in_295; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_295 <= _GEN_2436;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_296 <= io_rvfi_mem_data_in_296; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_296 <= _GEN_2437;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_297 <= io_rvfi_mem_data_in_297; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_297 <= _GEN_2438;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_298 <= io_rvfi_mem_data_in_298; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_298 <= _GEN_2439;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_299 <= io_rvfi_mem_data_in_299; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_299 <= _GEN_2440;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_300 <= io_rvfi_mem_data_in_300; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_300 <= _GEN_2441;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_301 <= io_rvfi_mem_data_in_301; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_301 <= _GEN_2442;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_302 <= io_rvfi_mem_data_in_302; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_302 <= _GEN_2443;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_303 <= io_rvfi_mem_data_in_303; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_303 <= _GEN_2444;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_304 <= io_rvfi_mem_data_in_304; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_304 <= _GEN_2445;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_305 <= io_rvfi_mem_data_in_305; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_305 <= _GEN_2446;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_306 <= io_rvfi_mem_data_in_306; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_306 <= _GEN_2447;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_307 <= io_rvfi_mem_data_in_307; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_307 <= _GEN_2448;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_308 <= io_rvfi_mem_data_in_308; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_308 <= _GEN_2449;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_309 <= io_rvfi_mem_data_in_309; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_309 <= _GEN_2450;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_310 <= io_rvfi_mem_data_in_310; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_310 <= _GEN_2451;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_311 <= io_rvfi_mem_data_in_311; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_311 <= _GEN_2452;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_312 <= io_rvfi_mem_data_in_312; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_312 <= _GEN_2453;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_313 <= io_rvfi_mem_data_in_313; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_313 <= _GEN_2454;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_314 <= io_rvfi_mem_data_in_314; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_314 <= _GEN_2455;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_315 <= io_rvfi_mem_data_in_315; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_315 <= _GEN_2456;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_316 <= io_rvfi_mem_data_in_316; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_316 <= _GEN_2457;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_317 <= io_rvfi_mem_data_in_317; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_317 <= _GEN_2458;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_318 <= io_rvfi_mem_data_in_318; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_318 <= _GEN_2459;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_319 <= io_rvfi_mem_data_in_319; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_319 <= _GEN_2460;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_320 <= io_rvfi_mem_data_in_320; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_320 <= _GEN_2461;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_321 <= io_rvfi_mem_data_in_321; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_321 <= _GEN_2462;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_322 <= io_rvfi_mem_data_in_322; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_322 <= _GEN_2463;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_323 <= io_rvfi_mem_data_in_323; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_323 <= _GEN_2464;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_324 <= io_rvfi_mem_data_in_324; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_324 <= _GEN_2465;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_325 <= io_rvfi_mem_data_in_325; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_325 <= _GEN_2466;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_326 <= io_rvfi_mem_data_in_326; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_326 <= _GEN_2467;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_327 <= io_rvfi_mem_data_in_327; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_327 <= _GEN_2468;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_328 <= io_rvfi_mem_data_in_328; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_328 <= _GEN_2469;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_329 <= io_rvfi_mem_data_in_329; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_329 <= _GEN_2470;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_330 <= io_rvfi_mem_data_in_330; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_330 <= _GEN_2471;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_331 <= io_rvfi_mem_data_in_331; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_331 <= _GEN_2472;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_332 <= io_rvfi_mem_data_in_332; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_332 <= _GEN_2473;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_333 <= io_rvfi_mem_data_in_333; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_333 <= _GEN_2474;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_334 <= io_rvfi_mem_data_in_334; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_334 <= _GEN_2475;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_335 <= io_rvfi_mem_data_in_335; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_335 <= _GEN_2476;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_336 <= io_rvfi_mem_data_in_336; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_336 <= _GEN_2477;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_337 <= io_rvfi_mem_data_in_337; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_337 <= _GEN_2478;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_338 <= io_rvfi_mem_data_in_338; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_338 <= _GEN_2479;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_339 <= io_rvfi_mem_data_in_339; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_339 <= _GEN_2480;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_340 <= io_rvfi_mem_data_in_340; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_340 <= _GEN_2481;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_341 <= io_rvfi_mem_data_in_341; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_341 <= _GEN_2482;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_342 <= io_rvfi_mem_data_in_342; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_342 <= _GEN_2483;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_343 <= io_rvfi_mem_data_in_343; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_343 <= _GEN_2484;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_344 <= io_rvfi_mem_data_in_344; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_344 <= _GEN_2485;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_345 <= io_rvfi_mem_data_in_345; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_345 <= _GEN_2486;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_346 <= io_rvfi_mem_data_in_346; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_346 <= _GEN_2487;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_347 <= io_rvfi_mem_data_in_347; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_347 <= _GEN_2488;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_348 <= io_rvfi_mem_data_in_348; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_348 <= _GEN_2489;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_349 <= io_rvfi_mem_data_in_349; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_349 <= _GEN_2490;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_350 <= io_rvfi_mem_data_in_350; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_350 <= _GEN_2491;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_351 <= io_rvfi_mem_data_in_351; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_351 <= _GEN_2492;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_352 <= io_rvfi_mem_data_in_352; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_352 <= _GEN_2493;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_353 <= io_rvfi_mem_data_in_353; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_353 <= _GEN_2494;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_354 <= io_rvfi_mem_data_in_354; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_354 <= _GEN_2495;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_355 <= io_rvfi_mem_data_in_355; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_355 <= _GEN_2496;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_356 <= io_rvfi_mem_data_in_356; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_356 <= _GEN_2497;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_357 <= io_rvfi_mem_data_in_357; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_357 <= _GEN_2498;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_358 <= io_rvfi_mem_data_in_358; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_358 <= _GEN_2499;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_359 <= io_rvfi_mem_data_in_359; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_359 <= _GEN_2500;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_360 <= io_rvfi_mem_data_in_360; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_360 <= _GEN_2501;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_361 <= io_rvfi_mem_data_in_361; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_361 <= _GEN_2502;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_362 <= io_rvfi_mem_data_in_362; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_362 <= _GEN_2503;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_363 <= io_rvfi_mem_data_in_363; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_363 <= _GEN_2504;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_364 <= io_rvfi_mem_data_in_364; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_364 <= _GEN_2505;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_365 <= io_rvfi_mem_data_in_365; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_365 <= _GEN_2506;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_366 <= io_rvfi_mem_data_in_366; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_366 <= _GEN_2507;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_367 <= io_rvfi_mem_data_in_367; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_367 <= _GEN_2508;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_368 <= io_rvfi_mem_data_in_368; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_368 <= _GEN_2509;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_369 <= io_rvfi_mem_data_in_369; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_369 <= _GEN_2510;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_370 <= io_rvfi_mem_data_in_370; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_370 <= _GEN_2511;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_371 <= io_rvfi_mem_data_in_371; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_371 <= _GEN_2512;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_372 <= io_rvfi_mem_data_in_372; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_372 <= _GEN_2513;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_373 <= io_rvfi_mem_data_in_373; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_373 <= _GEN_2514;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_374 <= io_rvfi_mem_data_in_374; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_374 <= _GEN_2515;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_375 <= io_rvfi_mem_data_in_375; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_375 <= _GEN_2516;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_376 <= io_rvfi_mem_data_in_376; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_376 <= _GEN_2517;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_377 <= io_rvfi_mem_data_in_377; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_377 <= _GEN_2518;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_378 <= io_rvfi_mem_data_in_378; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_378 <= _GEN_2519;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_379 <= io_rvfi_mem_data_in_379; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_379 <= _GEN_2520;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_380 <= io_rvfi_mem_data_in_380; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_380 <= _GEN_2521;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_381 <= io_rvfi_mem_data_in_381; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_381 <= _GEN_2522;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_382 <= io_rvfi_mem_data_in_382; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_382 <= _GEN_2523;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_383 <= io_rvfi_mem_data_in_383; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_383 <= _GEN_2524;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_384 <= io_rvfi_mem_data_in_384; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_384 <= _GEN_2525;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_385 <= io_rvfi_mem_data_in_385; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_385 <= _GEN_2526;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_386 <= io_rvfi_mem_data_in_386; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_386 <= _GEN_2527;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_387 <= io_rvfi_mem_data_in_387; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_387 <= _GEN_2528;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_388 <= io_rvfi_mem_data_in_388; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_388 <= _GEN_2529;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_389 <= io_rvfi_mem_data_in_389; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_389 <= _GEN_2530;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_390 <= io_rvfi_mem_data_in_390; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_390 <= _GEN_2531;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_391 <= io_rvfi_mem_data_in_391; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_391 <= _GEN_2532;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_392 <= io_rvfi_mem_data_in_392; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_392 <= _GEN_2533;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_393 <= io_rvfi_mem_data_in_393; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_393 <= _GEN_2534;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_394 <= io_rvfi_mem_data_in_394; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_394 <= _GEN_2535;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_395 <= io_rvfi_mem_data_in_395; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_395 <= _GEN_2536;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_396 <= io_rvfi_mem_data_in_396; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_396 <= _GEN_2537;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_397 <= io_rvfi_mem_data_in_397; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_397 <= _GEN_2538;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_398 <= io_rvfi_mem_data_in_398; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_398 <= _GEN_2539;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_399 <= io_rvfi_mem_data_in_399; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_399 <= _GEN_2540;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_400 <= io_rvfi_mem_data_in_400; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_400 <= _GEN_2541;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_401 <= io_rvfi_mem_data_in_401; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_401 <= _GEN_2542;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_402 <= io_rvfi_mem_data_in_402; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_402 <= _GEN_2543;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_403 <= io_rvfi_mem_data_in_403; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_403 <= _GEN_2544;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_404 <= io_rvfi_mem_data_in_404; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_404 <= _GEN_2545;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_405 <= io_rvfi_mem_data_in_405; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_405 <= _GEN_2546;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_406 <= io_rvfi_mem_data_in_406; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_406 <= _GEN_2547;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_407 <= io_rvfi_mem_data_in_407; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_407 <= _GEN_2548;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_408 <= io_rvfi_mem_data_in_408; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_408 <= _GEN_2549;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_409 <= io_rvfi_mem_data_in_409; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_409 <= _GEN_2550;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_410 <= io_rvfi_mem_data_in_410; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_410 <= _GEN_2551;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_411 <= io_rvfi_mem_data_in_411; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_411 <= _GEN_2552;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_412 <= io_rvfi_mem_data_in_412; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_412 <= _GEN_2553;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_413 <= io_rvfi_mem_data_in_413; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_413 <= _GEN_2554;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_414 <= io_rvfi_mem_data_in_414; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_414 <= _GEN_2555;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_415 <= io_rvfi_mem_data_in_415; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_415 <= _GEN_2556;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_416 <= io_rvfi_mem_data_in_416; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_416 <= _GEN_2557;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_417 <= io_rvfi_mem_data_in_417; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_417 <= _GEN_2558;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_418 <= io_rvfi_mem_data_in_418; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_418 <= _GEN_2559;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_419 <= io_rvfi_mem_data_in_419; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_419 <= _GEN_2560;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_420 <= io_rvfi_mem_data_in_420; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_420 <= _GEN_2561;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_421 <= io_rvfi_mem_data_in_421; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_421 <= _GEN_2562;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_422 <= io_rvfi_mem_data_in_422; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_422 <= _GEN_2563;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_423 <= io_rvfi_mem_data_in_423; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_423 <= _GEN_2564;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_424 <= io_rvfi_mem_data_in_424; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_424 <= _GEN_2565;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_425 <= io_rvfi_mem_data_in_425; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_425 <= _GEN_2566;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_426 <= io_rvfi_mem_data_in_426; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_426 <= _GEN_2567;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_427 <= io_rvfi_mem_data_in_427; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_427 <= _GEN_2568;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_428 <= io_rvfi_mem_data_in_428; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_428 <= _GEN_2569;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_429 <= io_rvfi_mem_data_in_429; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_429 <= _GEN_2570;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_430 <= io_rvfi_mem_data_in_430; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_430 <= _GEN_2571;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_431 <= io_rvfi_mem_data_in_431; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_431 <= _GEN_2572;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_432 <= io_rvfi_mem_data_in_432; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_432 <= _GEN_2573;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_433 <= io_rvfi_mem_data_in_433; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_433 <= _GEN_2574;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_434 <= io_rvfi_mem_data_in_434; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_434 <= _GEN_2575;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_435 <= io_rvfi_mem_data_in_435; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_435 <= _GEN_2576;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_436 <= io_rvfi_mem_data_in_436; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_436 <= _GEN_2577;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_437 <= io_rvfi_mem_data_in_437; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_437 <= _GEN_2578;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_438 <= io_rvfi_mem_data_in_438; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_438 <= _GEN_2579;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_439 <= io_rvfi_mem_data_in_439; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_439 <= _GEN_2580;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_440 <= io_rvfi_mem_data_in_440; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_440 <= _GEN_2581;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_441 <= io_rvfi_mem_data_in_441; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_441 <= _GEN_2582;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_442 <= io_rvfi_mem_data_in_442; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_442 <= _GEN_2583;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_443 <= io_rvfi_mem_data_in_443; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_443 <= _GEN_2584;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_444 <= io_rvfi_mem_data_in_444; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_444 <= _GEN_2585;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_445 <= io_rvfi_mem_data_in_445; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_445 <= _GEN_2586;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_446 <= io_rvfi_mem_data_in_446; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_446 <= _GEN_2587;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_447 <= io_rvfi_mem_data_in_447; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_447 <= _GEN_2588;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_448 <= io_rvfi_mem_data_in_448; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_448 <= _GEN_2589;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_449 <= io_rvfi_mem_data_in_449; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_449 <= _GEN_2590;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_450 <= io_rvfi_mem_data_in_450; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_450 <= _GEN_2591;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_451 <= io_rvfi_mem_data_in_451; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_451 <= _GEN_2592;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_452 <= io_rvfi_mem_data_in_452; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_452 <= _GEN_2593;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_453 <= io_rvfi_mem_data_in_453; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_453 <= _GEN_2594;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_454 <= io_rvfi_mem_data_in_454; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_454 <= _GEN_2595;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_455 <= io_rvfi_mem_data_in_455; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_455 <= _GEN_2596;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_456 <= io_rvfi_mem_data_in_456; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_456 <= _GEN_2597;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_457 <= io_rvfi_mem_data_in_457; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_457 <= _GEN_2598;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_458 <= io_rvfi_mem_data_in_458; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_458 <= _GEN_2599;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_459 <= io_rvfi_mem_data_in_459; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_459 <= _GEN_2600;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_460 <= io_rvfi_mem_data_in_460; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_460 <= _GEN_2601;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_461 <= io_rvfi_mem_data_in_461; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_461 <= _GEN_2602;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_462 <= io_rvfi_mem_data_in_462; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_462 <= _GEN_2603;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_463 <= io_rvfi_mem_data_in_463; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_463 <= _GEN_2604;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_464 <= io_rvfi_mem_data_in_464; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_464 <= _GEN_2605;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_465 <= io_rvfi_mem_data_in_465; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_465 <= _GEN_2606;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_466 <= io_rvfi_mem_data_in_466; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_466 <= _GEN_2607;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_467 <= io_rvfi_mem_data_in_467; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_467 <= _GEN_2608;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_468 <= io_rvfi_mem_data_in_468; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_468 <= _GEN_2609;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_469 <= io_rvfi_mem_data_in_469; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_469 <= _GEN_2610;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_470 <= io_rvfi_mem_data_in_470; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_470 <= _GEN_2611;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_471 <= io_rvfi_mem_data_in_471; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_471 <= _GEN_2612;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_472 <= io_rvfi_mem_data_in_472; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_472 <= _GEN_2613;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_473 <= io_rvfi_mem_data_in_473; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_473 <= _GEN_2614;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_474 <= io_rvfi_mem_data_in_474; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_474 <= _GEN_2615;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_475 <= io_rvfi_mem_data_in_475; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_475 <= _GEN_2616;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_476 <= io_rvfi_mem_data_in_476; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_476 <= _GEN_2617;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_477 <= io_rvfi_mem_data_in_477; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_477 <= _GEN_2618;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_478 <= io_rvfi_mem_data_in_478; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_478 <= _GEN_2619;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_479 <= io_rvfi_mem_data_in_479; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_479 <= _GEN_2620;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_480 <= io_rvfi_mem_data_in_480; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_480 <= _GEN_2621;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_481 <= io_rvfi_mem_data_in_481; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_481 <= _GEN_2622;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_482 <= io_rvfi_mem_data_in_482; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_482 <= _GEN_2623;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_483 <= io_rvfi_mem_data_in_483; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_483 <= _GEN_2624;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_484 <= io_rvfi_mem_data_in_484; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_484 <= _GEN_2625;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_485 <= io_rvfi_mem_data_in_485; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_485 <= _GEN_2626;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_486 <= io_rvfi_mem_data_in_486; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_486 <= _GEN_2627;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_487 <= io_rvfi_mem_data_in_487; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_487 <= _GEN_2628;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_488 <= io_rvfi_mem_data_in_488; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_488 <= _GEN_2629;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_489 <= io_rvfi_mem_data_in_489; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_489 <= _GEN_2630;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_490 <= io_rvfi_mem_data_in_490; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_490 <= _GEN_2631;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_491 <= io_rvfi_mem_data_in_491; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_491 <= _GEN_2632;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_492 <= io_rvfi_mem_data_in_492; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_492 <= _GEN_2633;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_493 <= io_rvfi_mem_data_in_493; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_493 <= _GEN_2634;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_494 <= io_rvfi_mem_data_in_494; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_494 <= _GEN_2635;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_495 <= io_rvfi_mem_data_in_495; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_495 <= _GEN_2636;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_496 <= io_rvfi_mem_data_in_496; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_496 <= _GEN_2637;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_497 <= io_rvfi_mem_data_in_497; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_497 <= _GEN_2638;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_498 <= io_rvfi_mem_data_in_498; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_498 <= _GEN_2639;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_499 <= io_rvfi_mem_data_in_499; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_499 <= _GEN_2640;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_500 <= io_rvfi_mem_data_in_500; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_500 <= _GEN_2641;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_501 <= io_rvfi_mem_data_in_501; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_501 <= _GEN_2642;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_502 <= io_rvfi_mem_data_in_502; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_502 <= _GEN_2643;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_503 <= io_rvfi_mem_data_in_503; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_503 <= _GEN_2644;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_504 <= io_rvfi_mem_data_in_504; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_504 <= _GEN_2645;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_505 <= io_rvfi_mem_data_in_505; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_505 <= _GEN_2646;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_506 <= io_rvfi_mem_data_in_506; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_506 <= _GEN_2647;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_507 <= io_rvfi_mem_data_in_507; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_507 <= _GEN_2648;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_508 <= io_rvfi_mem_data_in_508; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_508 <= _GEN_2649;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_509 <= io_rvfi_mem_data_in_509; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_509 <= _GEN_2650;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_510 <= io_rvfi_mem_data_in_510; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_510 <= _GEN_2651;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_511 <= io_rvfi_mem_data_in_511; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_511 <= _GEN_2652;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_512 <= io_rvfi_mem_data_in_512; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_512 <= _GEN_2653;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_513 <= io_rvfi_mem_data_in_513; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_513 <= _GEN_2654;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_514 <= io_rvfi_mem_data_in_514; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_514 <= _GEN_2655;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_515 <= io_rvfi_mem_data_in_515; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_515 <= _GEN_2656;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_516 <= io_rvfi_mem_data_in_516; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_516 <= _GEN_2657;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_517 <= io_rvfi_mem_data_in_517; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_517 <= _GEN_2658;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_518 <= io_rvfi_mem_data_in_518; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_518 <= _GEN_2659;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_519 <= io_rvfi_mem_data_in_519; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_519 <= _GEN_2660;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_520 <= io_rvfi_mem_data_in_520; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_520 <= _GEN_2661;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_521 <= io_rvfi_mem_data_in_521; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_521 <= _GEN_2662;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_522 <= io_rvfi_mem_data_in_522; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_522 <= _GEN_2663;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_523 <= io_rvfi_mem_data_in_523; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_523 <= _GEN_2664;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_524 <= io_rvfi_mem_data_in_524; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_524 <= _GEN_2665;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_525 <= io_rvfi_mem_data_in_525; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_525 <= _GEN_2666;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_526 <= io_rvfi_mem_data_in_526; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_526 <= _GEN_2667;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_527 <= io_rvfi_mem_data_in_527; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_527 <= _GEN_2668;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_528 <= io_rvfi_mem_data_in_528; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_528 <= _GEN_2669;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_529 <= io_rvfi_mem_data_in_529; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_529 <= _GEN_2670;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_530 <= io_rvfi_mem_data_in_530; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_530 <= _GEN_2671;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_531 <= io_rvfi_mem_data_in_531; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_531 <= _GEN_2672;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_532 <= io_rvfi_mem_data_in_532; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_532 <= _GEN_2673;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_533 <= io_rvfi_mem_data_in_533; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_533 <= _GEN_2674;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_534 <= io_rvfi_mem_data_in_534; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_534 <= _GEN_2675;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_535 <= io_rvfi_mem_data_in_535; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_535 <= _GEN_2676;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_536 <= io_rvfi_mem_data_in_536; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_536 <= _GEN_2677;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_537 <= io_rvfi_mem_data_in_537; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_537 <= _GEN_2678;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_538 <= io_rvfi_mem_data_in_538; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_538 <= _GEN_2679;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_539 <= io_rvfi_mem_data_in_539; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_539 <= _GEN_2680;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_540 <= io_rvfi_mem_data_in_540; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_540 <= _GEN_2681;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_541 <= io_rvfi_mem_data_in_541; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_541 <= _GEN_2682;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_542 <= io_rvfi_mem_data_in_542; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_542 <= _GEN_2683;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_543 <= io_rvfi_mem_data_in_543; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_543 <= _GEN_2684;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_544 <= io_rvfi_mem_data_in_544; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_544 <= _GEN_2685;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_545 <= io_rvfi_mem_data_in_545; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_545 <= _GEN_2686;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_546 <= io_rvfi_mem_data_in_546; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_546 <= _GEN_2687;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_547 <= io_rvfi_mem_data_in_547; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_547 <= _GEN_2688;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_548 <= io_rvfi_mem_data_in_548; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_548 <= _GEN_2689;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_549 <= io_rvfi_mem_data_in_549; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_549 <= _GEN_2690;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_550 <= io_rvfi_mem_data_in_550; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_550 <= _GEN_2691;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_551 <= io_rvfi_mem_data_in_551; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_551 <= _GEN_2692;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_552 <= io_rvfi_mem_data_in_552; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_552 <= _GEN_2693;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_553 <= io_rvfi_mem_data_in_553; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_553 <= _GEN_2694;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_554 <= io_rvfi_mem_data_in_554; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_554 <= _GEN_2695;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_555 <= io_rvfi_mem_data_in_555; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_555 <= _GEN_2696;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_556 <= io_rvfi_mem_data_in_556; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_556 <= _GEN_2697;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_557 <= io_rvfi_mem_data_in_557; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_557 <= _GEN_2698;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_558 <= io_rvfi_mem_data_in_558; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_558 <= _GEN_2699;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_559 <= io_rvfi_mem_data_in_559; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_559 <= _GEN_2700;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_560 <= io_rvfi_mem_data_in_560; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_560 <= _GEN_2701;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_561 <= io_rvfi_mem_data_in_561; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_561 <= _GEN_2702;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_562 <= io_rvfi_mem_data_in_562; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_562 <= _GEN_2703;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_563 <= io_rvfi_mem_data_in_563; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_563 <= _GEN_2704;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_564 <= io_rvfi_mem_data_in_564; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_564 <= _GEN_2705;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_565 <= io_rvfi_mem_data_in_565; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_565 <= _GEN_2706;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_566 <= io_rvfi_mem_data_in_566; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_566 <= _GEN_2707;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_567 <= io_rvfi_mem_data_in_567; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_567 <= _GEN_2708;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_568 <= io_rvfi_mem_data_in_568; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_568 <= _GEN_2709;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_569 <= io_rvfi_mem_data_in_569; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_569 <= _GEN_2710;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_570 <= io_rvfi_mem_data_in_570; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_570 <= _GEN_2711;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_571 <= io_rvfi_mem_data_in_571; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_571 <= _GEN_2712;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_572 <= io_rvfi_mem_data_in_572; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_572 <= _GEN_2713;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_573 <= io_rvfi_mem_data_in_573; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_573 <= _GEN_2714;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_574 <= io_rvfi_mem_data_in_574; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_574 <= _GEN_2715;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_575 <= io_rvfi_mem_data_in_575; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_575 <= _GEN_2716;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_576 <= io_rvfi_mem_data_in_576; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_576 <= _GEN_2717;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_577 <= io_rvfi_mem_data_in_577; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_577 <= _GEN_2718;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_578 <= io_rvfi_mem_data_in_578; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_578 <= _GEN_2719;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_579 <= io_rvfi_mem_data_in_579; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_579 <= _GEN_2720;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_580 <= io_rvfi_mem_data_in_580; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_580 <= _GEN_2721;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_581 <= io_rvfi_mem_data_in_581; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_581 <= _GEN_2722;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_582 <= io_rvfi_mem_data_in_582; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_582 <= _GEN_2723;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_583 <= io_rvfi_mem_data_in_583; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_583 <= _GEN_2724;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_584 <= io_rvfi_mem_data_in_584; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_584 <= _GEN_2725;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_585 <= io_rvfi_mem_data_in_585; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_585 <= _GEN_2726;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_586 <= io_rvfi_mem_data_in_586; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_586 <= _GEN_2727;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_587 <= io_rvfi_mem_data_in_587; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_587 <= _GEN_2728;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_588 <= io_rvfi_mem_data_in_588; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_588 <= _GEN_2729;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_589 <= io_rvfi_mem_data_in_589; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_589 <= _GEN_2730;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_590 <= io_rvfi_mem_data_in_590; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_590 <= _GEN_2731;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_591 <= io_rvfi_mem_data_in_591; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_591 <= _GEN_2732;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_592 <= io_rvfi_mem_data_in_592; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_592 <= _GEN_2733;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_593 <= io_rvfi_mem_data_in_593; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_593 <= _GEN_2734;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_594 <= io_rvfi_mem_data_in_594; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_594 <= _GEN_2735;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_595 <= io_rvfi_mem_data_in_595; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_595 <= _GEN_2736;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_596 <= io_rvfi_mem_data_in_596; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_596 <= _GEN_2737;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_597 <= io_rvfi_mem_data_in_597; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_597 <= _GEN_2738;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_598 <= io_rvfi_mem_data_in_598; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_598 <= _GEN_2739;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_599 <= io_rvfi_mem_data_in_599; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_599 <= _GEN_2740;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_600 <= io_rvfi_mem_data_in_600; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_600 <= _GEN_2741;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_601 <= io_rvfi_mem_data_in_601; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_601 <= _GEN_2742;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_602 <= io_rvfi_mem_data_in_602; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_602 <= _GEN_2743;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_603 <= io_rvfi_mem_data_in_603; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_603 <= _GEN_2744;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_604 <= io_rvfi_mem_data_in_604; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_604 <= _GEN_2745;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_605 <= io_rvfi_mem_data_in_605; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_605 <= _GEN_2746;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_606 <= io_rvfi_mem_data_in_606; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_606 <= _GEN_2747;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_607 <= io_rvfi_mem_data_in_607; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_607 <= _GEN_2748;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_608 <= io_rvfi_mem_data_in_608; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_608 <= _GEN_2749;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_609 <= io_rvfi_mem_data_in_609; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_609 <= _GEN_2750;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_610 <= io_rvfi_mem_data_in_610; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_610 <= _GEN_2751;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_611 <= io_rvfi_mem_data_in_611; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_611 <= _GEN_2752;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_612 <= io_rvfi_mem_data_in_612; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_612 <= _GEN_2753;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_613 <= io_rvfi_mem_data_in_613; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_613 <= _GEN_2754;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_614 <= io_rvfi_mem_data_in_614; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_614 <= _GEN_2755;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_615 <= io_rvfi_mem_data_in_615; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_615 <= _GEN_2756;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_616 <= io_rvfi_mem_data_in_616; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_616 <= _GEN_2757;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_617 <= io_rvfi_mem_data_in_617; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_617 <= _GEN_2758;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_618 <= io_rvfi_mem_data_in_618; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_618 <= _GEN_2759;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_619 <= io_rvfi_mem_data_in_619; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_619 <= _GEN_2760;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_620 <= io_rvfi_mem_data_in_620; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_620 <= _GEN_2761;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_621 <= io_rvfi_mem_data_in_621; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_621 <= _GEN_2762;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_622 <= io_rvfi_mem_data_in_622; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_622 <= _GEN_2763;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_623 <= io_rvfi_mem_data_in_623; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_623 <= _GEN_2764;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_624 <= io_rvfi_mem_data_in_624; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_624 <= _GEN_2765;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_625 <= io_rvfi_mem_data_in_625; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_625 <= _GEN_2766;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_626 <= io_rvfi_mem_data_in_626; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_626 <= _GEN_2767;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_627 <= io_rvfi_mem_data_in_627; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_627 <= _GEN_2768;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_628 <= io_rvfi_mem_data_in_628; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_628 <= _GEN_2769;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_629 <= io_rvfi_mem_data_in_629; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_629 <= _GEN_2770;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_630 <= io_rvfi_mem_data_in_630; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_630 <= _GEN_2771;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_631 <= io_rvfi_mem_data_in_631; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_631 <= _GEN_2772;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_632 <= io_rvfi_mem_data_in_632; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_632 <= _GEN_2773;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_633 <= io_rvfi_mem_data_in_633; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_633 <= _GEN_2774;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_634 <= io_rvfi_mem_data_in_634; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_634 <= _GEN_2775;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_635 <= io_rvfi_mem_data_in_635; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_635 <= _GEN_2776;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_636 <= io_rvfi_mem_data_in_636; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_636 <= _GEN_2777;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_637 <= io_rvfi_mem_data_in_637; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_637 <= _GEN_2778;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_638 <= io_rvfi_mem_data_in_638; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_638 <= _GEN_2779;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_639 <= io_rvfi_mem_data_in_639; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_639 <= _GEN_2780;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_640 <= io_rvfi_mem_data_in_640; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_640 <= _GEN_2781;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_641 <= io_rvfi_mem_data_in_641; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_641 <= _GEN_2782;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_642 <= io_rvfi_mem_data_in_642; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_642 <= _GEN_2783;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_643 <= io_rvfi_mem_data_in_643; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_643 <= _GEN_2784;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_644 <= io_rvfi_mem_data_in_644; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_644 <= _GEN_2785;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_645 <= io_rvfi_mem_data_in_645; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_645 <= _GEN_2786;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_646 <= io_rvfi_mem_data_in_646; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_646 <= _GEN_2787;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_647 <= io_rvfi_mem_data_in_647; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_647 <= _GEN_2788;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_648 <= io_rvfi_mem_data_in_648; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_648 <= _GEN_2789;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_649 <= io_rvfi_mem_data_in_649; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_649 <= _GEN_2790;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_650 <= io_rvfi_mem_data_in_650; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_650 <= _GEN_2791;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_651 <= io_rvfi_mem_data_in_651; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_651 <= _GEN_2792;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_652 <= io_rvfi_mem_data_in_652; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_652 <= _GEN_2793;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_653 <= io_rvfi_mem_data_in_653; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_653 <= _GEN_2794;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_654 <= io_rvfi_mem_data_in_654; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_654 <= _GEN_2795;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_655 <= io_rvfi_mem_data_in_655; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_655 <= _GEN_2796;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_656 <= io_rvfi_mem_data_in_656; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_656 <= _GEN_2797;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_657 <= io_rvfi_mem_data_in_657; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_657 <= _GEN_2798;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_658 <= io_rvfi_mem_data_in_658; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_658 <= _GEN_2799;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_659 <= io_rvfi_mem_data_in_659; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_659 <= _GEN_2800;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_660 <= io_rvfi_mem_data_in_660; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_660 <= _GEN_2801;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_661 <= io_rvfi_mem_data_in_661; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_661 <= _GEN_2802;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_662 <= io_rvfi_mem_data_in_662; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_662 <= _GEN_2803;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_663 <= io_rvfi_mem_data_in_663; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_663 <= _GEN_2804;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_664 <= io_rvfi_mem_data_in_664; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_664 <= _GEN_2805;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_665 <= io_rvfi_mem_data_in_665; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_665 <= _GEN_2806;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_666 <= io_rvfi_mem_data_in_666; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_666 <= _GEN_2807;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_667 <= io_rvfi_mem_data_in_667; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_667 <= _GEN_2808;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_668 <= io_rvfi_mem_data_in_668; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_668 <= _GEN_2809;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_669 <= io_rvfi_mem_data_in_669; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_669 <= _GEN_2810;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_670 <= io_rvfi_mem_data_in_670; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_670 <= _GEN_2811;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_671 <= io_rvfi_mem_data_in_671; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_671 <= _GEN_2812;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_672 <= io_rvfi_mem_data_in_672; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_672 <= _GEN_2813;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_673 <= io_rvfi_mem_data_in_673; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_673 <= _GEN_2814;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_674 <= io_rvfi_mem_data_in_674; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_674 <= _GEN_2815;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_675 <= io_rvfi_mem_data_in_675; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_675 <= _GEN_2816;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_676 <= io_rvfi_mem_data_in_676; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_676 <= _GEN_2817;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_677 <= io_rvfi_mem_data_in_677; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_677 <= _GEN_2818;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_678 <= io_rvfi_mem_data_in_678; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_678 <= _GEN_2819;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_679 <= io_rvfi_mem_data_in_679; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_679 <= _GEN_2820;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_680 <= io_rvfi_mem_data_in_680; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_680 <= _GEN_2821;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_681 <= io_rvfi_mem_data_in_681; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_681 <= _GEN_2822;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_682 <= io_rvfi_mem_data_in_682; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_682 <= _GEN_2823;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_683 <= io_rvfi_mem_data_in_683; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_683 <= _GEN_2824;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_684 <= io_rvfi_mem_data_in_684; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_684 <= _GEN_2825;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_685 <= io_rvfi_mem_data_in_685; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_685 <= _GEN_2826;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_686 <= io_rvfi_mem_data_in_686; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_686 <= _GEN_2827;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_687 <= io_rvfi_mem_data_in_687; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_687 <= _GEN_2828;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_688 <= io_rvfi_mem_data_in_688; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_688 <= _GEN_2829;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_689 <= io_rvfi_mem_data_in_689; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_689 <= _GEN_2830;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_690 <= io_rvfi_mem_data_in_690; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_690 <= _GEN_2831;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_691 <= io_rvfi_mem_data_in_691; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_691 <= _GEN_2832;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_692 <= io_rvfi_mem_data_in_692; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_692 <= _GEN_2833;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_693 <= io_rvfi_mem_data_in_693; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_693 <= _GEN_2834;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_694 <= io_rvfi_mem_data_in_694; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_694 <= _GEN_2835;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_695 <= io_rvfi_mem_data_in_695; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_695 <= _GEN_2836;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_696 <= io_rvfi_mem_data_in_696; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_696 <= _GEN_2837;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_697 <= io_rvfi_mem_data_in_697; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_697 <= _GEN_2838;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_698 <= io_rvfi_mem_data_in_698; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_698 <= _GEN_2839;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_699 <= io_rvfi_mem_data_in_699; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_699 <= _GEN_2840;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_700 <= io_rvfi_mem_data_in_700; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_700 <= _GEN_2841;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_701 <= io_rvfi_mem_data_in_701; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_701 <= _GEN_2842;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_702 <= io_rvfi_mem_data_in_702; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_702 <= _GEN_2843;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_703 <= io_rvfi_mem_data_in_703; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_703 <= _GEN_2844;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_704 <= io_rvfi_mem_data_in_704; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_704 <= _GEN_2845;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_705 <= io_rvfi_mem_data_in_705; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_705 <= _GEN_2846;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_706 <= io_rvfi_mem_data_in_706; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_706 <= _GEN_2847;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_707 <= io_rvfi_mem_data_in_707; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_707 <= _GEN_2848;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_708 <= io_rvfi_mem_data_in_708; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_708 <= _GEN_2849;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_709 <= io_rvfi_mem_data_in_709; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_709 <= _GEN_2850;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_710 <= io_rvfi_mem_data_in_710; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_710 <= _GEN_2851;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_711 <= io_rvfi_mem_data_in_711; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_711 <= _GEN_2852;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_712 <= io_rvfi_mem_data_in_712; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_712 <= _GEN_2853;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_713 <= io_rvfi_mem_data_in_713; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_713 <= _GEN_2854;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_714 <= io_rvfi_mem_data_in_714; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_714 <= _GEN_2855;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_715 <= io_rvfi_mem_data_in_715; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_715 <= _GEN_2856;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_716 <= io_rvfi_mem_data_in_716; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_716 <= _GEN_2857;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_717 <= io_rvfi_mem_data_in_717; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_717 <= _GEN_2858;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_718 <= io_rvfi_mem_data_in_718; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_718 <= _GEN_2859;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_719 <= io_rvfi_mem_data_in_719; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_719 <= _GEN_2860;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_720 <= io_rvfi_mem_data_in_720; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_720 <= _GEN_2861;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_721 <= io_rvfi_mem_data_in_721; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_721 <= _GEN_2862;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_722 <= io_rvfi_mem_data_in_722; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_722 <= _GEN_2863;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_723 <= io_rvfi_mem_data_in_723; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_723 <= _GEN_2864;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_724 <= io_rvfi_mem_data_in_724; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_724 <= _GEN_2865;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_725 <= io_rvfi_mem_data_in_725; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_725 <= _GEN_2866;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_726 <= io_rvfi_mem_data_in_726; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_726 <= _GEN_2867;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_727 <= io_rvfi_mem_data_in_727; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_727 <= _GEN_2868;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_728 <= io_rvfi_mem_data_in_728; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_728 <= _GEN_2869;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_729 <= io_rvfi_mem_data_in_729; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_729 <= _GEN_2870;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_730 <= io_rvfi_mem_data_in_730; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_730 <= _GEN_2871;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_731 <= io_rvfi_mem_data_in_731; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_731 <= _GEN_2872;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_732 <= io_rvfi_mem_data_in_732; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_732 <= _GEN_2873;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_733 <= io_rvfi_mem_data_in_733; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_733 <= _GEN_2874;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_734 <= io_rvfi_mem_data_in_734; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_734 <= _GEN_2875;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_735 <= io_rvfi_mem_data_in_735; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_735 <= _GEN_2876;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_736 <= io_rvfi_mem_data_in_736; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_736 <= _GEN_2877;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_737 <= io_rvfi_mem_data_in_737; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_737 <= _GEN_2878;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_738 <= io_rvfi_mem_data_in_738; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_738 <= _GEN_2879;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_739 <= io_rvfi_mem_data_in_739; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_739 <= _GEN_2880;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_740 <= io_rvfi_mem_data_in_740; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_740 <= _GEN_2881;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_741 <= io_rvfi_mem_data_in_741; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_741 <= _GEN_2882;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_742 <= io_rvfi_mem_data_in_742; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_742 <= _GEN_2883;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_743 <= io_rvfi_mem_data_in_743; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_743 <= _GEN_2884;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_744 <= io_rvfi_mem_data_in_744; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_744 <= _GEN_2885;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_745 <= io_rvfi_mem_data_in_745; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_745 <= _GEN_2886;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_746 <= io_rvfi_mem_data_in_746; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_746 <= _GEN_2887;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_747 <= io_rvfi_mem_data_in_747; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_747 <= _GEN_2888;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_748 <= io_rvfi_mem_data_in_748; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_748 <= _GEN_2889;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_749 <= io_rvfi_mem_data_in_749; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_749 <= _GEN_2890;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_750 <= io_rvfi_mem_data_in_750; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_750 <= _GEN_2891;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_751 <= io_rvfi_mem_data_in_751; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_751 <= _GEN_2892;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_752 <= io_rvfi_mem_data_in_752; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_752 <= _GEN_2893;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_753 <= io_rvfi_mem_data_in_753; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_753 <= _GEN_2894;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_754 <= io_rvfi_mem_data_in_754; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_754 <= _GEN_2895;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_755 <= io_rvfi_mem_data_in_755; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_755 <= _GEN_2896;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_756 <= io_rvfi_mem_data_in_756; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_756 <= _GEN_2897;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_757 <= io_rvfi_mem_data_in_757; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_757 <= _GEN_2898;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_758 <= io_rvfi_mem_data_in_758; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_758 <= _GEN_2899;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_759 <= io_rvfi_mem_data_in_759; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_759 <= _GEN_2900;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_760 <= io_rvfi_mem_data_in_760; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_760 <= _GEN_2901;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_761 <= io_rvfi_mem_data_in_761; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_761 <= _GEN_2902;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_762 <= io_rvfi_mem_data_in_762; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_762 <= _GEN_2903;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_763 <= io_rvfi_mem_data_in_763; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_763 <= _GEN_2904;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_764 <= io_rvfi_mem_data_in_764; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_764 <= _GEN_2905;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_765 <= io_rvfi_mem_data_in_765; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_765 <= _GEN_2906;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_766 <= io_rvfi_mem_data_in_766; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_766 <= _GEN_2907;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_767 <= io_rvfi_mem_data_in_767; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_767 <= _GEN_2908;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_768 <= io_rvfi_mem_data_in_768; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_768 <= _GEN_2909;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_769 <= io_rvfi_mem_data_in_769; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_769 <= _GEN_2910;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_770 <= io_rvfi_mem_data_in_770; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_770 <= _GEN_2911;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_771 <= io_rvfi_mem_data_in_771; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_771 <= _GEN_2912;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_772 <= io_rvfi_mem_data_in_772; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_772 <= _GEN_2913;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_773 <= io_rvfi_mem_data_in_773; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_773 <= _GEN_2914;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_774 <= io_rvfi_mem_data_in_774; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_774 <= _GEN_2915;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_775 <= io_rvfi_mem_data_in_775; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_775 <= _GEN_2916;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_776 <= io_rvfi_mem_data_in_776; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_776 <= _GEN_2917;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_777 <= io_rvfi_mem_data_in_777; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_777 <= _GEN_2918;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_778 <= io_rvfi_mem_data_in_778; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_778 <= _GEN_2919;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_779 <= io_rvfi_mem_data_in_779; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_779 <= _GEN_2920;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_780 <= io_rvfi_mem_data_in_780; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_780 <= _GEN_2921;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_781 <= io_rvfi_mem_data_in_781; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_781 <= _GEN_2922;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_782 <= io_rvfi_mem_data_in_782; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_782 <= _GEN_2923;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_783 <= io_rvfi_mem_data_in_783; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_783 <= _GEN_2924;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_784 <= io_rvfi_mem_data_in_784; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_784 <= _GEN_2925;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_785 <= io_rvfi_mem_data_in_785; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_785 <= _GEN_2926;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_786 <= io_rvfi_mem_data_in_786; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_786 <= _GEN_2927;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_787 <= io_rvfi_mem_data_in_787; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_787 <= _GEN_2928;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_788 <= io_rvfi_mem_data_in_788; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_788 <= _GEN_2929;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_789 <= io_rvfi_mem_data_in_789; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_789 <= _GEN_2930;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_790 <= io_rvfi_mem_data_in_790; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_790 <= _GEN_2931;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_791 <= io_rvfi_mem_data_in_791; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_791 <= _GEN_2932;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_792 <= io_rvfi_mem_data_in_792; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_792 <= _GEN_2933;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_793 <= io_rvfi_mem_data_in_793; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_793 <= _GEN_2934;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_794 <= io_rvfi_mem_data_in_794; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_794 <= _GEN_2935;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_795 <= io_rvfi_mem_data_in_795; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_795 <= _GEN_2936;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_796 <= io_rvfi_mem_data_in_796; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_796 <= _GEN_2937;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_797 <= io_rvfi_mem_data_in_797; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_797 <= _GEN_2938;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_798 <= io_rvfi_mem_data_in_798; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_798 <= _GEN_2939;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_799 <= io_rvfi_mem_data_in_799; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_799 <= _GEN_2940;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_800 <= io_rvfi_mem_data_in_800; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_800 <= _GEN_2941;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_801 <= io_rvfi_mem_data_in_801; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_801 <= _GEN_2942;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_802 <= io_rvfi_mem_data_in_802; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_802 <= _GEN_2943;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_803 <= io_rvfi_mem_data_in_803; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_803 <= _GEN_2944;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_804 <= io_rvfi_mem_data_in_804; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_804 <= _GEN_2945;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_805 <= io_rvfi_mem_data_in_805; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_805 <= _GEN_2946;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_806 <= io_rvfi_mem_data_in_806; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_806 <= _GEN_2947;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_807 <= io_rvfi_mem_data_in_807; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_807 <= _GEN_2948;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_808 <= io_rvfi_mem_data_in_808; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_808 <= _GEN_2949;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_809 <= io_rvfi_mem_data_in_809; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_809 <= _GEN_2950;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_810 <= io_rvfi_mem_data_in_810; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_810 <= _GEN_2951;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_811 <= io_rvfi_mem_data_in_811; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_811 <= _GEN_2952;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_812 <= io_rvfi_mem_data_in_812; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_812 <= _GEN_2953;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_813 <= io_rvfi_mem_data_in_813; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_813 <= _GEN_2954;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_814 <= io_rvfi_mem_data_in_814; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_814 <= _GEN_2955;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_815 <= io_rvfi_mem_data_in_815; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_815 <= _GEN_2956;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_816 <= io_rvfi_mem_data_in_816; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_816 <= _GEN_2957;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_817 <= io_rvfi_mem_data_in_817; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_817 <= _GEN_2958;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_818 <= io_rvfi_mem_data_in_818; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_818 <= _GEN_2959;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_819 <= io_rvfi_mem_data_in_819; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_819 <= _GEN_2960;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_820 <= io_rvfi_mem_data_in_820; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_820 <= _GEN_2961;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_821 <= io_rvfi_mem_data_in_821; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_821 <= _GEN_2962;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_822 <= io_rvfi_mem_data_in_822; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_822 <= _GEN_2963;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_823 <= io_rvfi_mem_data_in_823; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_823 <= _GEN_2964;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_824 <= io_rvfi_mem_data_in_824; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_824 <= _GEN_2965;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_825 <= io_rvfi_mem_data_in_825; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_825 <= _GEN_2966;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_826 <= io_rvfi_mem_data_in_826; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_826 <= _GEN_2967;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_827 <= io_rvfi_mem_data_in_827; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_827 <= _GEN_2968;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_828 <= io_rvfi_mem_data_in_828; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_828 <= _GEN_2969;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_829 <= io_rvfi_mem_data_in_829; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_829 <= _GEN_2970;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_830 <= io_rvfi_mem_data_in_830; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_830 <= _GEN_2971;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_831 <= io_rvfi_mem_data_in_831; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_831 <= _GEN_2972;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_832 <= io_rvfi_mem_data_in_832; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_832 <= _GEN_2973;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_833 <= io_rvfi_mem_data_in_833; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_833 <= _GEN_2974;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_834 <= io_rvfi_mem_data_in_834; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_834 <= _GEN_2975;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_835 <= io_rvfi_mem_data_in_835; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_835 <= _GEN_2976;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_836 <= io_rvfi_mem_data_in_836; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_836 <= _GEN_2977;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_837 <= io_rvfi_mem_data_in_837; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_837 <= _GEN_2978;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_838 <= io_rvfi_mem_data_in_838; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_838 <= _GEN_2979;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_839 <= io_rvfi_mem_data_in_839; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_839 <= _GEN_2980;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_840 <= io_rvfi_mem_data_in_840; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_840 <= _GEN_2981;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_841 <= io_rvfi_mem_data_in_841; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_841 <= _GEN_2982;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_842 <= io_rvfi_mem_data_in_842; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_842 <= _GEN_2983;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_843 <= io_rvfi_mem_data_in_843; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_843 <= _GEN_2984;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_844 <= io_rvfi_mem_data_in_844; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_844 <= _GEN_2985;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_845 <= io_rvfi_mem_data_in_845; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_845 <= _GEN_2986;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_846 <= io_rvfi_mem_data_in_846; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_846 <= _GEN_2987;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_847 <= io_rvfi_mem_data_in_847; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_847 <= _GEN_2988;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_848 <= io_rvfi_mem_data_in_848; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_848 <= _GEN_2989;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_849 <= io_rvfi_mem_data_in_849; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_849 <= _GEN_2990;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_850 <= io_rvfi_mem_data_in_850; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_850 <= _GEN_2991;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_851 <= io_rvfi_mem_data_in_851; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_851 <= _GEN_2992;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_852 <= io_rvfi_mem_data_in_852; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_852 <= _GEN_2993;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_853 <= io_rvfi_mem_data_in_853; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_853 <= _GEN_2994;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_854 <= io_rvfi_mem_data_in_854; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_854 <= _GEN_2995;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_855 <= io_rvfi_mem_data_in_855; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_855 <= _GEN_2996;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_856 <= io_rvfi_mem_data_in_856; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_856 <= _GEN_2997;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_857 <= io_rvfi_mem_data_in_857; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_857 <= _GEN_2998;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_858 <= io_rvfi_mem_data_in_858; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_858 <= _GEN_2999;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_859 <= io_rvfi_mem_data_in_859; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_859 <= _GEN_3000;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_860 <= io_rvfi_mem_data_in_860; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_860 <= _GEN_3001;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_861 <= io_rvfi_mem_data_in_861; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_861 <= _GEN_3002;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_862 <= io_rvfi_mem_data_in_862; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_862 <= _GEN_3003;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_863 <= io_rvfi_mem_data_in_863; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_863 <= _GEN_3004;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_864 <= io_rvfi_mem_data_in_864; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_864 <= _GEN_3005;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_865 <= io_rvfi_mem_data_in_865; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_865 <= _GEN_3006;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_866 <= io_rvfi_mem_data_in_866; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_866 <= _GEN_3007;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_867 <= io_rvfi_mem_data_in_867; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_867 <= _GEN_3008;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_868 <= io_rvfi_mem_data_in_868; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_868 <= _GEN_3009;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_869 <= io_rvfi_mem_data_in_869; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_869 <= _GEN_3010;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_870 <= io_rvfi_mem_data_in_870; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_870 <= _GEN_3011;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_871 <= io_rvfi_mem_data_in_871; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_871 <= _GEN_3012;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_872 <= io_rvfi_mem_data_in_872; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_872 <= _GEN_3013;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_873 <= io_rvfi_mem_data_in_873; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_873 <= _GEN_3014;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_874 <= io_rvfi_mem_data_in_874; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_874 <= _GEN_3015;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_875 <= io_rvfi_mem_data_in_875; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_875 <= _GEN_3016;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_876 <= io_rvfi_mem_data_in_876; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_876 <= _GEN_3017;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_877 <= io_rvfi_mem_data_in_877; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_877 <= _GEN_3018;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_878 <= io_rvfi_mem_data_in_878; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_878 <= _GEN_3019;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_879 <= io_rvfi_mem_data_in_879; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_879 <= _GEN_3020;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_880 <= io_rvfi_mem_data_in_880; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_880 <= _GEN_3021;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_881 <= io_rvfi_mem_data_in_881; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_881 <= _GEN_3022;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_882 <= io_rvfi_mem_data_in_882; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_882 <= _GEN_3023;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_883 <= io_rvfi_mem_data_in_883; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_883 <= _GEN_3024;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_884 <= io_rvfi_mem_data_in_884; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_884 <= _GEN_3025;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_885 <= io_rvfi_mem_data_in_885; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_885 <= _GEN_3026;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_886 <= io_rvfi_mem_data_in_886; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_886 <= _GEN_3027;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_887 <= io_rvfi_mem_data_in_887; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_887 <= _GEN_3028;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_888 <= io_rvfi_mem_data_in_888; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_888 <= _GEN_3029;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_889 <= io_rvfi_mem_data_in_889; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_889 <= _GEN_3030;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_890 <= io_rvfi_mem_data_in_890; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_890 <= _GEN_3031;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_891 <= io_rvfi_mem_data_in_891; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_891 <= _GEN_3032;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_892 <= io_rvfi_mem_data_in_892; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_892 <= _GEN_3033;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_893 <= io_rvfi_mem_data_in_893; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_893 <= _GEN_3034;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_894 <= io_rvfi_mem_data_in_894; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_894 <= _GEN_3035;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_895 <= io_rvfi_mem_data_in_895; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_895 <= _GEN_3036;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_896 <= io_rvfi_mem_data_in_896; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_896 <= _GEN_3037;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_897 <= io_rvfi_mem_data_in_897; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_897 <= _GEN_3038;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_898 <= io_rvfi_mem_data_in_898; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_898 <= _GEN_3039;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_899 <= io_rvfi_mem_data_in_899; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_899 <= _GEN_3040;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_900 <= io_rvfi_mem_data_in_900; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_900 <= _GEN_3041;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_901 <= io_rvfi_mem_data_in_901; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_901 <= _GEN_3042;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_902 <= io_rvfi_mem_data_in_902; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_902 <= _GEN_3043;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_903 <= io_rvfi_mem_data_in_903; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_903 <= _GEN_3044;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_904 <= io_rvfi_mem_data_in_904; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_904 <= _GEN_3045;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_905 <= io_rvfi_mem_data_in_905; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_905 <= _GEN_3046;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_906 <= io_rvfi_mem_data_in_906; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_906 <= _GEN_3047;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_907 <= io_rvfi_mem_data_in_907; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_907 <= _GEN_3048;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_908 <= io_rvfi_mem_data_in_908; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_908 <= _GEN_3049;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_909 <= io_rvfi_mem_data_in_909; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_909 <= _GEN_3050;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_910 <= io_rvfi_mem_data_in_910; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_910 <= _GEN_3051;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_911 <= io_rvfi_mem_data_in_911; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_911 <= _GEN_3052;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_912 <= io_rvfi_mem_data_in_912; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_912 <= _GEN_3053;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_913 <= io_rvfi_mem_data_in_913; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_913 <= _GEN_3054;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_914 <= io_rvfi_mem_data_in_914; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_914 <= _GEN_3055;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_915 <= io_rvfi_mem_data_in_915; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_915 <= _GEN_3056;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_916 <= io_rvfi_mem_data_in_916; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_916 <= _GEN_3057;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_917 <= io_rvfi_mem_data_in_917; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_917 <= _GEN_3058;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_918 <= io_rvfi_mem_data_in_918; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_918 <= _GEN_3059;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_919 <= io_rvfi_mem_data_in_919; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_919 <= _GEN_3060;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_920 <= io_rvfi_mem_data_in_920; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_920 <= _GEN_3061;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_921 <= io_rvfi_mem_data_in_921; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_921 <= _GEN_3062;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_922 <= io_rvfi_mem_data_in_922; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_922 <= _GEN_3063;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_923 <= io_rvfi_mem_data_in_923; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_923 <= _GEN_3064;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_924 <= io_rvfi_mem_data_in_924; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_924 <= _GEN_3065;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_925 <= io_rvfi_mem_data_in_925; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_925 <= _GEN_3066;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_926 <= io_rvfi_mem_data_in_926; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_926 <= _GEN_3067;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_927 <= io_rvfi_mem_data_in_927; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_927 <= _GEN_3068;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_928 <= io_rvfi_mem_data_in_928; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_928 <= _GEN_3069;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_929 <= io_rvfi_mem_data_in_929; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_929 <= _GEN_3070;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_930 <= io_rvfi_mem_data_in_930; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_930 <= _GEN_3071;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_931 <= io_rvfi_mem_data_in_931; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_931 <= _GEN_3072;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_932 <= io_rvfi_mem_data_in_932; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_932 <= _GEN_3073;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_933 <= io_rvfi_mem_data_in_933; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_933 <= _GEN_3074;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_934 <= io_rvfi_mem_data_in_934; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_934 <= _GEN_3075;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_935 <= io_rvfi_mem_data_in_935; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_935 <= _GEN_3076;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_936 <= io_rvfi_mem_data_in_936; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_936 <= _GEN_3077;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_937 <= io_rvfi_mem_data_in_937; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_937 <= _GEN_3078;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_938 <= io_rvfi_mem_data_in_938; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_938 <= _GEN_3079;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_939 <= io_rvfi_mem_data_in_939; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_939 <= _GEN_3080;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_940 <= io_rvfi_mem_data_in_940; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_940 <= _GEN_3081;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_941 <= io_rvfi_mem_data_in_941; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_941 <= _GEN_3082;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_942 <= io_rvfi_mem_data_in_942; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_942 <= _GEN_3083;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_943 <= io_rvfi_mem_data_in_943; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_943 <= _GEN_3084;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_944 <= io_rvfi_mem_data_in_944; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_944 <= _GEN_3085;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_945 <= io_rvfi_mem_data_in_945; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_945 <= _GEN_3086;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_946 <= io_rvfi_mem_data_in_946; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_946 <= _GEN_3087;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_947 <= io_rvfi_mem_data_in_947; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_947 <= _GEN_3088;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_948 <= io_rvfi_mem_data_in_948; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_948 <= _GEN_3089;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_949 <= io_rvfi_mem_data_in_949; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_949 <= _GEN_3090;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_950 <= io_rvfi_mem_data_in_950; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_950 <= _GEN_3091;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_951 <= io_rvfi_mem_data_in_951; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_951 <= _GEN_3092;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_952 <= io_rvfi_mem_data_in_952; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_952 <= _GEN_3093;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_953 <= io_rvfi_mem_data_in_953; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_953 <= _GEN_3094;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_954 <= io_rvfi_mem_data_in_954; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_954 <= _GEN_3095;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_955 <= io_rvfi_mem_data_in_955; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_955 <= _GEN_3096;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_956 <= io_rvfi_mem_data_in_956; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_956 <= _GEN_3097;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_957 <= io_rvfi_mem_data_in_957; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_957 <= _GEN_3098;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_958 <= io_rvfi_mem_data_in_958; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_958 <= _GEN_3099;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_959 <= io_rvfi_mem_data_in_959; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_959 <= _GEN_3100;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_960 <= io_rvfi_mem_data_in_960; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_960 <= _GEN_3101;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_961 <= io_rvfi_mem_data_in_961; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_961 <= _GEN_3102;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_962 <= io_rvfi_mem_data_in_962; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_962 <= _GEN_3103;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_963 <= io_rvfi_mem_data_in_963; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_963 <= _GEN_3104;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_964 <= io_rvfi_mem_data_in_964; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_964 <= _GEN_3105;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_965 <= io_rvfi_mem_data_in_965; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_965 <= _GEN_3106;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_966 <= io_rvfi_mem_data_in_966; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_966 <= _GEN_3107;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_967 <= io_rvfi_mem_data_in_967; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_967 <= _GEN_3108;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_968 <= io_rvfi_mem_data_in_968; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_968 <= _GEN_3109;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_969 <= io_rvfi_mem_data_in_969; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_969 <= _GEN_3110;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_970 <= io_rvfi_mem_data_in_970; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_970 <= _GEN_3111;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_971 <= io_rvfi_mem_data_in_971; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_971 <= _GEN_3112;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_972 <= io_rvfi_mem_data_in_972; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_972 <= _GEN_3113;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_973 <= io_rvfi_mem_data_in_973; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_973 <= _GEN_3114;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_974 <= io_rvfi_mem_data_in_974; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_974 <= _GEN_3115;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_975 <= io_rvfi_mem_data_in_975; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_975 <= _GEN_3116;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_976 <= io_rvfi_mem_data_in_976; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_976 <= _GEN_3117;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_977 <= io_rvfi_mem_data_in_977; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_977 <= _GEN_3118;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_978 <= io_rvfi_mem_data_in_978; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_978 <= _GEN_3119;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_979 <= io_rvfi_mem_data_in_979; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_979 <= _GEN_3120;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_980 <= io_rvfi_mem_data_in_980; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_980 <= _GEN_3121;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_981 <= io_rvfi_mem_data_in_981; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_981 <= _GEN_3122;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_982 <= io_rvfi_mem_data_in_982; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_982 <= _GEN_3123;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_983 <= io_rvfi_mem_data_in_983; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_983 <= _GEN_3124;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_984 <= io_rvfi_mem_data_in_984; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_984 <= _GEN_3125;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_985 <= io_rvfi_mem_data_in_985; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_985 <= _GEN_3126;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_986 <= io_rvfi_mem_data_in_986; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_986 <= _GEN_3127;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_987 <= io_rvfi_mem_data_in_987; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_987 <= _GEN_3128;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_988 <= io_rvfi_mem_data_in_988; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_988 <= _GEN_3129;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_989 <= io_rvfi_mem_data_in_989; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_989 <= _GEN_3130;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_990 <= io_rvfi_mem_data_in_990; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_990 <= _GEN_3131;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_991 <= io_rvfi_mem_data_in_991; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_991 <= _GEN_3132;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_992 <= io_rvfi_mem_data_in_992; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_992 <= _GEN_3133;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_993 <= io_rvfi_mem_data_in_993; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_993 <= _GEN_3134;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_994 <= io_rvfi_mem_data_in_994; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_994 <= _GEN_3135;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_995 <= io_rvfi_mem_data_in_995; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_995 <= _GEN_3136;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_996 <= io_rvfi_mem_data_in_996; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_996 <= _GEN_3137;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_997 <= io_rvfi_mem_data_in_997; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_997 <= _GEN_3138;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_998 <= io_rvfi_mem_data_in_998; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_998 <= _GEN_3139;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_999 <= io_rvfi_mem_data_in_999; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_999 <= _GEN_3140;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1000 <= io_rvfi_mem_data_in_1000; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1000 <= _GEN_3141;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1001 <= io_rvfi_mem_data_in_1001; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1001 <= _GEN_3142;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1002 <= io_rvfi_mem_data_in_1002; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1002 <= _GEN_3143;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1003 <= io_rvfi_mem_data_in_1003; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1003 <= _GEN_3144;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1004 <= io_rvfi_mem_data_in_1004; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1004 <= _GEN_3145;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1005 <= io_rvfi_mem_data_in_1005; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1005 <= _GEN_3146;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1006 <= io_rvfi_mem_data_in_1006; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1006 <= _GEN_3147;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1007 <= io_rvfi_mem_data_in_1007; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1007 <= _GEN_3148;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1008 <= io_rvfi_mem_data_in_1008; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1008 <= _GEN_3149;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1009 <= io_rvfi_mem_data_in_1009; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1009 <= _GEN_3150;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1010 <= io_rvfi_mem_data_in_1010; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1010 <= _GEN_3151;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1011 <= io_rvfi_mem_data_in_1011; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1011 <= _GEN_3152;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1012 <= io_rvfi_mem_data_in_1012; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1012 <= _GEN_3153;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1013 <= io_rvfi_mem_data_in_1013; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1013 <= _GEN_3154;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1014 <= io_rvfi_mem_data_in_1014; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1014 <= _GEN_3155;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1015 <= io_rvfi_mem_data_in_1015; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1015 <= _GEN_3156;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1016 <= io_rvfi_mem_data_in_1016; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1016 <= _GEN_3157;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1017 <= io_rvfi_mem_data_in_1017; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1017 <= _GEN_3158;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1018 <= io_rvfi_mem_data_in_1018; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1018 <= _GEN_3159;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1019 <= io_rvfi_mem_data_in_1019; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1019 <= _GEN_3160;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1020 <= io_rvfi_mem_data_in_1020; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1020 <= _GEN_3161;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1021 <= io_rvfi_mem_data_in_1021; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1021 <= _GEN_3162;
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      DMemory_1022 <= io_rvfi_mem_data_in_1022; // @[cpu.scala 71:17]
    end else if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
      if (!(_stall_T)) begin // @[cpu.scala 198:32]
        if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
          DMemory_1022 <= _GEN_3163;
        end
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 196:29]
        if (!(_stall_T)) begin // @[cpu.scala 198:32]
          if (EXMEMop == 7'h23) begin // @[cpu.scala 200:32]
            DMemory_1023 <= _GEN_3164;
          end
        end
      end
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      IMemory_0 <= io_rvfi_insn_in_0; // @[cpu.scala 65:18]
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      IMemory_1 <= io_rvfi_insn_in_1; // @[cpu.scala 65:18]
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      IMemory_2 <= io_rvfi_insn_in_2; // @[cpu.scala 65:18]
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      IMemory_3 <= io_rvfi_insn_in_3; // @[cpu.scala 65:18]
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      IMemory_4 <= io_rvfi_insn_in_4; // @[cpu.scala 65:18]
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      IMemory_5 <= io_rvfi_insn_in_5; // @[cpu.scala 65:18]
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      IMemory_6 <= io_rvfi_insn_in_6; // @[cpu.scala 65:18]
    end
    if (io_rvfi_rst) begin // @[cpu.scala 55:21]
      IMemory_7 <= io_rvfi_insn_in_7; // @[cpu.scala 65:18]
    end
    if (reset) begin // @[cpu.scala 48:49]
      IFIDIR <= 32'h13; // @[cpu.scala 48:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      if (~stall) begin // @[cpu.scala 117:27]
        if (~takeBranch) begin // @[cpu.scala 118:34]
          IFIDIR <= _GEN_1023; // @[cpu.scala 121:16]
        end else begin
          IFIDIR <= 32'h13; // @[cpu.scala 125:16]
        end
      end
    end
    if (reset) begin // @[cpu.scala 48:49]
      IDEXIR <= 32'h13; // @[cpu.scala 48:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      if (~stall) begin // @[cpu.scala 117:27]
        IDEXIR <= IFIDIR; // @[cpu.scala 170:14]
      end else begin
        IDEXIR <= 32'h13; // @[cpu.scala 172:14]
      end
    end
    if (reset) begin // @[cpu.scala 48:49]
      EXMEMIR <= 32'h13; // @[cpu.scala 48:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      EXMEMIR <= IDEXIR; // @[cpu.scala 192:13]
    end
    if (reset) begin // @[cpu.scala 48:49]
      MEMWBIR <= 32'h13; // @[cpu.scala 48:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      MEMWBIR <= EXMEMIR; // @[cpu.scala 204:13]
    end
    if (reset) begin // @[cpu.scala 51:22]
      CurPC <= 64'h0; // @[cpu.scala 51:22]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 55:21]
      if (~stall) begin // @[cpu.scala 117:27]
        CurPC <= PC; // @[cpu.scala 141:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  PC = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  Regs_0 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  Regs_1 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  Regs_2 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  Regs_3 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  Regs_4 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  Regs_5 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  Regs_6 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  Regs_7 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  Regs_8 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  Regs_9 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  Regs_10 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  Regs_11 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  Regs_12 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  Regs_13 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  Regs_14 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  Regs_15 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  Regs_16 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  Regs_17 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  Regs_18 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  Regs_19 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  Regs_20 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  Regs_21 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  Regs_22 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  Regs_23 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  Regs_24 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  Regs_25 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  Regs_26 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  Regs_27 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  Regs_28 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  Regs_29 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  Regs_30 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  Regs_31 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  IDEXA = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  IDEXB = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  EXMEMB = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  EXMEMALUOut = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  MEMWBValue = _RAND_37[63:0];
  _RAND_38 = {1{`RANDOM}};
  DMemory_0 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  DMemory_1 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  DMemory_2 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  DMemory_3 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  DMemory_4 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  DMemory_5 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  DMemory_6 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  DMemory_7 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  DMemory_8 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  DMemory_9 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  DMemory_10 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  DMemory_11 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  DMemory_12 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  DMemory_13 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  DMemory_14 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  DMemory_15 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  DMemory_16 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  DMemory_17 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  DMemory_18 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  DMemory_19 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  DMemory_20 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  DMemory_21 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  DMemory_22 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  DMemory_23 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  DMemory_24 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  DMemory_25 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  DMemory_26 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  DMemory_27 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  DMemory_28 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  DMemory_29 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  DMemory_30 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  DMemory_31 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  DMemory_32 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  DMemory_33 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  DMemory_34 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  DMemory_35 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  DMemory_36 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  DMemory_37 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  DMemory_38 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  DMemory_39 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  DMemory_40 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  DMemory_41 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  DMemory_42 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  DMemory_43 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  DMemory_44 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  DMemory_45 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  DMemory_46 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  DMemory_47 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  DMemory_48 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  DMemory_49 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  DMemory_50 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  DMemory_51 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  DMemory_52 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  DMemory_53 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  DMemory_54 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  DMemory_55 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  DMemory_56 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  DMemory_57 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  DMemory_58 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  DMemory_59 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  DMemory_60 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  DMemory_61 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  DMemory_62 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  DMemory_63 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  DMemory_64 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  DMemory_65 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  DMemory_66 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  DMemory_67 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  DMemory_68 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  DMemory_69 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  DMemory_70 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  DMemory_71 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  DMemory_72 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  DMemory_73 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  DMemory_74 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  DMemory_75 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  DMemory_76 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  DMemory_77 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  DMemory_78 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  DMemory_79 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  DMemory_80 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  DMemory_81 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  DMemory_82 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  DMemory_83 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  DMemory_84 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  DMemory_85 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  DMemory_86 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  DMemory_87 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  DMemory_88 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  DMemory_89 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  DMemory_90 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  DMemory_91 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  DMemory_92 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  DMemory_93 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  DMemory_94 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  DMemory_95 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  DMemory_96 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  DMemory_97 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  DMemory_98 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  DMemory_99 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  DMemory_100 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  DMemory_101 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  DMemory_102 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  DMemory_103 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  DMemory_104 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  DMemory_105 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  DMemory_106 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  DMemory_107 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  DMemory_108 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  DMemory_109 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  DMemory_110 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  DMemory_111 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  DMemory_112 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  DMemory_113 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  DMemory_114 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  DMemory_115 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  DMemory_116 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  DMemory_117 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  DMemory_118 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  DMemory_119 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  DMemory_120 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  DMemory_121 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  DMemory_122 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  DMemory_123 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  DMemory_124 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  DMemory_125 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  DMemory_126 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  DMemory_127 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  DMemory_128 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  DMemory_129 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  DMemory_130 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  DMemory_131 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  DMemory_132 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  DMemory_133 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  DMemory_134 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  DMemory_135 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  DMemory_136 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  DMemory_137 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  DMemory_138 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  DMemory_139 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  DMemory_140 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  DMemory_141 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  DMemory_142 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  DMemory_143 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  DMemory_144 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  DMemory_145 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  DMemory_146 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  DMemory_147 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  DMemory_148 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  DMemory_149 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  DMemory_150 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  DMemory_151 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  DMemory_152 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  DMemory_153 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  DMemory_154 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  DMemory_155 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  DMemory_156 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  DMemory_157 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  DMemory_158 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  DMemory_159 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  DMemory_160 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  DMemory_161 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  DMemory_162 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  DMemory_163 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  DMemory_164 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  DMemory_165 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  DMemory_166 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  DMemory_167 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  DMemory_168 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  DMemory_169 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  DMemory_170 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  DMemory_171 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  DMemory_172 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  DMemory_173 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  DMemory_174 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  DMemory_175 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  DMemory_176 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  DMemory_177 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  DMemory_178 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  DMemory_179 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  DMemory_180 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  DMemory_181 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  DMemory_182 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  DMemory_183 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  DMemory_184 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  DMemory_185 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  DMemory_186 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  DMemory_187 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  DMemory_188 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  DMemory_189 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  DMemory_190 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  DMemory_191 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  DMemory_192 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  DMemory_193 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  DMemory_194 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  DMemory_195 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  DMemory_196 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  DMemory_197 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  DMemory_198 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  DMemory_199 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  DMemory_200 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  DMemory_201 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  DMemory_202 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  DMemory_203 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  DMemory_204 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  DMemory_205 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  DMemory_206 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  DMemory_207 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  DMemory_208 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  DMemory_209 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  DMemory_210 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  DMemory_211 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  DMemory_212 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  DMemory_213 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  DMemory_214 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  DMemory_215 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  DMemory_216 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  DMemory_217 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  DMemory_218 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  DMemory_219 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  DMemory_220 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  DMemory_221 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  DMemory_222 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  DMemory_223 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  DMemory_224 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  DMemory_225 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  DMemory_226 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  DMemory_227 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  DMemory_228 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  DMemory_229 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  DMemory_230 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  DMemory_231 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  DMemory_232 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  DMemory_233 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  DMemory_234 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  DMemory_235 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  DMemory_236 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  DMemory_237 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  DMemory_238 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  DMemory_239 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  DMemory_240 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  DMemory_241 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  DMemory_242 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  DMemory_243 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  DMemory_244 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  DMemory_245 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  DMemory_246 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  DMemory_247 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  DMemory_248 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  DMemory_249 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  DMemory_250 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  DMemory_251 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  DMemory_252 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  DMemory_253 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  DMemory_254 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  DMemory_255 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  DMemory_256 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  DMemory_257 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  DMemory_258 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  DMemory_259 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  DMemory_260 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  DMemory_261 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  DMemory_262 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  DMemory_263 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  DMemory_264 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  DMemory_265 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  DMemory_266 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  DMemory_267 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  DMemory_268 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  DMemory_269 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  DMemory_270 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  DMemory_271 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  DMemory_272 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  DMemory_273 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  DMemory_274 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  DMemory_275 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  DMemory_276 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  DMemory_277 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  DMemory_278 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  DMemory_279 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  DMemory_280 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  DMemory_281 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  DMemory_282 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  DMemory_283 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  DMemory_284 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  DMemory_285 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  DMemory_286 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  DMemory_287 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  DMemory_288 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  DMemory_289 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  DMemory_290 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  DMemory_291 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  DMemory_292 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  DMemory_293 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  DMemory_294 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  DMemory_295 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  DMemory_296 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  DMemory_297 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  DMemory_298 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  DMemory_299 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  DMemory_300 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  DMemory_301 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  DMemory_302 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  DMemory_303 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  DMemory_304 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  DMemory_305 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  DMemory_306 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  DMemory_307 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  DMemory_308 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  DMemory_309 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  DMemory_310 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  DMemory_311 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  DMemory_312 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  DMemory_313 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  DMemory_314 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  DMemory_315 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  DMemory_316 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  DMemory_317 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  DMemory_318 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  DMemory_319 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  DMemory_320 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  DMemory_321 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  DMemory_322 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  DMemory_323 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  DMemory_324 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  DMemory_325 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  DMemory_326 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  DMemory_327 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  DMemory_328 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  DMemory_329 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  DMemory_330 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  DMemory_331 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  DMemory_332 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  DMemory_333 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  DMemory_334 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  DMemory_335 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  DMemory_336 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  DMemory_337 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  DMemory_338 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  DMemory_339 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  DMemory_340 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  DMemory_341 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  DMemory_342 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  DMemory_343 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  DMemory_344 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  DMemory_345 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  DMemory_346 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  DMemory_347 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  DMemory_348 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  DMemory_349 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  DMemory_350 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  DMemory_351 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  DMemory_352 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  DMemory_353 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  DMemory_354 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  DMemory_355 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  DMemory_356 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  DMemory_357 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  DMemory_358 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  DMemory_359 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  DMemory_360 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  DMemory_361 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  DMemory_362 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  DMemory_363 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  DMemory_364 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  DMemory_365 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  DMemory_366 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  DMemory_367 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  DMemory_368 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  DMemory_369 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  DMemory_370 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  DMemory_371 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  DMemory_372 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  DMemory_373 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  DMemory_374 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  DMemory_375 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  DMemory_376 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  DMemory_377 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  DMemory_378 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  DMemory_379 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  DMemory_380 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  DMemory_381 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  DMemory_382 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  DMemory_383 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  DMemory_384 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  DMemory_385 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  DMemory_386 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  DMemory_387 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  DMemory_388 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  DMemory_389 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  DMemory_390 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  DMemory_391 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  DMemory_392 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  DMemory_393 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  DMemory_394 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  DMemory_395 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  DMemory_396 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  DMemory_397 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  DMemory_398 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  DMemory_399 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  DMemory_400 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  DMemory_401 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  DMemory_402 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  DMemory_403 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  DMemory_404 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  DMemory_405 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  DMemory_406 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  DMemory_407 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  DMemory_408 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  DMemory_409 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  DMemory_410 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  DMemory_411 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  DMemory_412 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  DMemory_413 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  DMemory_414 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  DMemory_415 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  DMemory_416 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  DMemory_417 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  DMemory_418 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  DMemory_419 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  DMemory_420 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  DMemory_421 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  DMemory_422 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  DMemory_423 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  DMemory_424 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  DMemory_425 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  DMemory_426 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  DMemory_427 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  DMemory_428 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  DMemory_429 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  DMemory_430 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  DMemory_431 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  DMemory_432 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  DMemory_433 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  DMemory_434 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  DMemory_435 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  DMemory_436 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  DMemory_437 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  DMemory_438 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  DMemory_439 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  DMemory_440 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  DMemory_441 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  DMemory_442 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  DMemory_443 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  DMemory_444 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  DMemory_445 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  DMemory_446 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  DMemory_447 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  DMemory_448 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  DMemory_449 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  DMemory_450 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  DMemory_451 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  DMemory_452 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  DMemory_453 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  DMemory_454 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  DMemory_455 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  DMemory_456 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  DMemory_457 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  DMemory_458 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  DMemory_459 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  DMemory_460 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  DMemory_461 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  DMemory_462 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  DMemory_463 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  DMemory_464 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  DMemory_465 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  DMemory_466 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  DMemory_467 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  DMemory_468 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  DMemory_469 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  DMemory_470 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  DMemory_471 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  DMemory_472 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  DMemory_473 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  DMemory_474 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  DMemory_475 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  DMemory_476 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  DMemory_477 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  DMemory_478 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  DMemory_479 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  DMemory_480 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  DMemory_481 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  DMemory_482 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  DMemory_483 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  DMemory_484 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  DMemory_485 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  DMemory_486 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  DMemory_487 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  DMemory_488 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  DMemory_489 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  DMemory_490 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  DMemory_491 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  DMemory_492 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  DMemory_493 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  DMemory_494 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  DMemory_495 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  DMemory_496 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  DMemory_497 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  DMemory_498 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  DMemory_499 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  DMemory_500 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  DMemory_501 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  DMemory_502 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  DMemory_503 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  DMemory_504 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  DMemory_505 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  DMemory_506 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  DMemory_507 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  DMemory_508 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  DMemory_509 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  DMemory_510 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  DMemory_511 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  DMemory_512 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  DMemory_513 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  DMemory_514 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  DMemory_515 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  DMemory_516 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  DMemory_517 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  DMemory_518 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  DMemory_519 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  DMemory_520 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  DMemory_521 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  DMemory_522 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  DMemory_523 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  DMemory_524 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  DMemory_525 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  DMemory_526 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  DMemory_527 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  DMemory_528 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  DMemory_529 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  DMemory_530 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  DMemory_531 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  DMemory_532 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  DMemory_533 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  DMemory_534 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  DMemory_535 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  DMemory_536 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  DMemory_537 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  DMemory_538 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  DMemory_539 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  DMemory_540 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  DMemory_541 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  DMemory_542 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  DMemory_543 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  DMemory_544 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  DMemory_545 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  DMemory_546 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  DMemory_547 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  DMemory_548 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  DMemory_549 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  DMemory_550 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  DMemory_551 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  DMemory_552 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  DMemory_553 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  DMemory_554 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  DMemory_555 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  DMemory_556 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  DMemory_557 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  DMemory_558 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  DMemory_559 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  DMemory_560 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  DMemory_561 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  DMemory_562 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  DMemory_563 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  DMemory_564 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  DMemory_565 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  DMemory_566 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  DMemory_567 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  DMemory_568 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  DMemory_569 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  DMemory_570 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  DMemory_571 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  DMemory_572 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  DMemory_573 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  DMemory_574 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  DMemory_575 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  DMemory_576 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  DMemory_577 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  DMemory_578 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  DMemory_579 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  DMemory_580 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  DMemory_581 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  DMemory_582 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  DMemory_583 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  DMemory_584 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  DMemory_585 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  DMemory_586 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  DMemory_587 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  DMemory_588 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  DMemory_589 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  DMemory_590 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  DMemory_591 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  DMemory_592 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  DMemory_593 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  DMemory_594 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  DMemory_595 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  DMemory_596 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  DMemory_597 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  DMemory_598 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  DMemory_599 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  DMemory_600 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  DMemory_601 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  DMemory_602 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  DMemory_603 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  DMemory_604 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  DMemory_605 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  DMemory_606 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  DMemory_607 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  DMemory_608 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  DMemory_609 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  DMemory_610 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  DMemory_611 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  DMemory_612 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  DMemory_613 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  DMemory_614 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  DMemory_615 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  DMemory_616 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  DMemory_617 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  DMemory_618 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  DMemory_619 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  DMemory_620 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  DMemory_621 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  DMemory_622 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  DMemory_623 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  DMemory_624 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  DMemory_625 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  DMemory_626 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  DMemory_627 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  DMemory_628 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  DMemory_629 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  DMemory_630 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  DMemory_631 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  DMemory_632 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  DMemory_633 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  DMemory_634 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  DMemory_635 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  DMemory_636 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  DMemory_637 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  DMemory_638 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  DMemory_639 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  DMemory_640 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  DMemory_641 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  DMemory_642 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  DMemory_643 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  DMemory_644 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  DMemory_645 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  DMemory_646 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  DMemory_647 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  DMemory_648 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  DMemory_649 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  DMemory_650 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  DMemory_651 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  DMemory_652 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  DMemory_653 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  DMemory_654 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  DMemory_655 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  DMemory_656 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  DMemory_657 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  DMemory_658 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  DMemory_659 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  DMemory_660 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  DMemory_661 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  DMemory_662 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  DMemory_663 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  DMemory_664 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  DMemory_665 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  DMemory_666 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  DMemory_667 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  DMemory_668 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  DMemory_669 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  DMemory_670 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  DMemory_671 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  DMemory_672 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  DMemory_673 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  DMemory_674 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  DMemory_675 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  DMemory_676 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  DMemory_677 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  DMemory_678 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  DMemory_679 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  DMemory_680 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  DMemory_681 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  DMemory_682 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  DMemory_683 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  DMemory_684 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  DMemory_685 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  DMemory_686 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  DMemory_687 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  DMemory_688 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  DMemory_689 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  DMemory_690 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  DMemory_691 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  DMemory_692 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  DMemory_693 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  DMemory_694 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  DMemory_695 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  DMemory_696 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  DMemory_697 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  DMemory_698 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  DMemory_699 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  DMemory_700 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  DMemory_701 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  DMemory_702 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  DMemory_703 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  DMemory_704 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  DMemory_705 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  DMemory_706 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  DMemory_707 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  DMemory_708 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  DMemory_709 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  DMemory_710 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  DMemory_711 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  DMemory_712 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  DMemory_713 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  DMemory_714 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  DMemory_715 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  DMemory_716 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  DMemory_717 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  DMemory_718 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  DMemory_719 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  DMemory_720 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  DMemory_721 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  DMemory_722 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  DMemory_723 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  DMemory_724 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  DMemory_725 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  DMemory_726 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  DMemory_727 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  DMemory_728 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  DMemory_729 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  DMemory_730 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  DMemory_731 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  DMemory_732 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  DMemory_733 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  DMemory_734 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  DMemory_735 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  DMemory_736 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  DMemory_737 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  DMemory_738 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  DMemory_739 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  DMemory_740 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  DMemory_741 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  DMemory_742 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  DMemory_743 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  DMemory_744 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  DMemory_745 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  DMemory_746 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  DMemory_747 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  DMemory_748 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  DMemory_749 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  DMemory_750 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  DMemory_751 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  DMemory_752 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  DMemory_753 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  DMemory_754 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  DMemory_755 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  DMemory_756 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  DMemory_757 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  DMemory_758 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  DMemory_759 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  DMemory_760 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  DMemory_761 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  DMemory_762 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  DMemory_763 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  DMemory_764 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  DMemory_765 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  DMemory_766 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  DMemory_767 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  DMemory_768 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  DMemory_769 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  DMemory_770 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  DMemory_771 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  DMemory_772 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  DMemory_773 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  DMemory_774 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  DMemory_775 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  DMemory_776 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  DMemory_777 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  DMemory_778 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  DMemory_779 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  DMemory_780 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  DMemory_781 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  DMemory_782 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  DMemory_783 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  DMemory_784 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  DMemory_785 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  DMemory_786 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  DMemory_787 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  DMemory_788 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  DMemory_789 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  DMemory_790 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  DMemory_791 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  DMemory_792 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  DMemory_793 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  DMemory_794 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  DMemory_795 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  DMemory_796 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  DMemory_797 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  DMemory_798 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  DMemory_799 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  DMemory_800 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  DMemory_801 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  DMemory_802 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  DMemory_803 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  DMemory_804 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  DMemory_805 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  DMemory_806 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  DMemory_807 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  DMemory_808 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  DMemory_809 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  DMemory_810 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  DMemory_811 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  DMemory_812 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  DMemory_813 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  DMemory_814 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  DMemory_815 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  DMemory_816 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  DMemory_817 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  DMemory_818 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  DMemory_819 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  DMemory_820 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  DMemory_821 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  DMemory_822 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  DMemory_823 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  DMemory_824 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  DMemory_825 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  DMemory_826 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  DMemory_827 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  DMemory_828 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  DMemory_829 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  DMemory_830 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  DMemory_831 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  DMemory_832 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  DMemory_833 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  DMemory_834 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  DMemory_835 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  DMemory_836 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  DMemory_837 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  DMemory_838 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  DMemory_839 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  DMemory_840 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  DMemory_841 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  DMemory_842 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  DMemory_843 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  DMemory_844 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  DMemory_845 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  DMemory_846 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  DMemory_847 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  DMemory_848 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  DMemory_849 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  DMemory_850 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  DMemory_851 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  DMemory_852 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  DMemory_853 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  DMemory_854 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  DMemory_855 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  DMemory_856 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  DMemory_857 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  DMemory_858 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  DMemory_859 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  DMemory_860 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  DMemory_861 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  DMemory_862 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  DMemory_863 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  DMemory_864 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  DMemory_865 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  DMemory_866 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  DMemory_867 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  DMemory_868 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  DMemory_869 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  DMemory_870 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  DMemory_871 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  DMemory_872 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  DMemory_873 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  DMemory_874 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  DMemory_875 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  DMemory_876 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  DMemory_877 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  DMemory_878 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  DMemory_879 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  DMemory_880 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  DMemory_881 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  DMemory_882 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  DMemory_883 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  DMemory_884 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  DMemory_885 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  DMemory_886 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  DMemory_887 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  DMemory_888 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  DMemory_889 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  DMemory_890 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  DMemory_891 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  DMemory_892 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  DMemory_893 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  DMemory_894 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  DMemory_895 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  DMemory_896 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  DMemory_897 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  DMemory_898 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  DMemory_899 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  DMemory_900 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  DMemory_901 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  DMemory_902 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  DMemory_903 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  DMemory_904 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  DMemory_905 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  DMemory_906 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  DMemory_907 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  DMemory_908 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  DMemory_909 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  DMemory_910 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  DMemory_911 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  DMemory_912 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  DMemory_913 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  DMemory_914 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  DMemory_915 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  DMemory_916 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  DMemory_917 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  DMemory_918 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  DMemory_919 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  DMemory_920 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  DMemory_921 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  DMemory_922 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  DMemory_923 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  DMemory_924 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  DMemory_925 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  DMemory_926 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  DMemory_927 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  DMemory_928 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  DMemory_929 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  DMemory_930 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  DMemory_931 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  DMemory_932 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  DMemory_933 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  DMemory_934 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  DMemory_935 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  DMemory_936 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  DMemory_937 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  DMemory_938 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  DMemory_939 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  DMemory_940 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  DMemory_941 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  DMemory_942 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  DMemory_943 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  DMemory_944 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  DMemory_945 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  DMemory_946 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  DMemory_947 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  DMemory_948 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  DMemory_949 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  DMemory_950 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  DMemory_951 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  DMemory_952 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  DMemory_953 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  DMemory_954 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  DMemory_955 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  DMemory_956 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  DMemory_957 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  DMemory_958 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  DMemory_959 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  DMemory_960 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  DMemory_961 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  DMemory_962 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  DMemory_963 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  DMemory_964 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  DMemory_965 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  DMemory_966 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  DMemory_967 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  DMemory_968 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  DMemory_969 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  DMemory_970 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  DMemory_971 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  DMemory_972 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  DMemory_973 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  DMemory_974 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  DMemory_975 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  DMemory_976 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  DMemory_977 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  DMemory_978 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  DMemory_979 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  DMemory_980 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  DMemory_981 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  DMemory_982 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  DMemory_983 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  DMemory_984 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  DMemory_985 = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  DMemory_986 = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  DMemory_987 = _RAND_1025[31:0];
  _RAND_1026 = {1{`RANDOM}};
  DMemory_988 = _RAND_1026[31:0];
  _RAND_1027 = {1{`RANDOM}};
  DMemory_989 = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  DMemory_990 = _RAND_1028[31:0];
  _RAND_1029 = {1{`RANDOM}};
  DMemory_991 = _RAND_1029[31:0];
  _RAND_1030 = {1{`RANDOM}};
  DMemory_992 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  DMemory_993 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  DMemory_994 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  DMemory_995 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  DMemory_996 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  DMemory_997 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  DMemory_998 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  DMemory_999 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  DMemory_1000 = _RAND_1038[31:0];
  _RAND_1039 = {1{`RANDOM}};
  DMemory_1001 = _RAND_1039[31:0];
  _RAND_1040 = {1{`RANDOM}};
  DMemory_1002 = _RAND_1040[31:0];
  _RAND_1041 = {1{`RANDOM}};
  DMemory_1003 = _RAND_1041[31:0];
  _RAND_1042 = {1{`RANDOM}};
  DMemory_1004 = _RAND_1042[31:0];
  _RAND_1043 = {1{`RANDOM}};
  DMemory_1005 = _RAND_1043[31:0];
  _RAND_1044 = {1{`RANDOM}};
  DMemory_1006 = _RAND_1044[31:0];
  _RAND_1045 = {1{`RANDOM}};
  DMemory_1007 = _RAND_1045[31:0];
  _RAND_1046 = {1{`RANDOM}};
  DMemory_1008 = _RAND_1046[31:0];
  _RAND_1047 = {1{`RANDOM}};
  DMemory_1009 = _RAND_1047[31:0];
  _RAND_1048 = {1{`RANDOM}};
  DMemory_1010 = _RAND_1048[31:0];
  _RAND_1049 = {1{`RANDOM}};
  DMemory_1011 = _RAND_1049[31:0];
  _RAND_1050 = {1{`RANDOM}};
  DMemory_1012 = _RAND_1050[31:0];
  _RAND_1051 = {1{`RANDOM}};
  DMemory_1013 = _RAND_1051[31:0];
  _RAND_1052 = {1{`RANDOM}};
  DMemory_1014 = _RAND_1052[31:0];
  _RAND_1053 = {1{`RANDOM}};
  DMemory_1015 = _RAND_1053[31:0];
  _RAND_1054 = {1{`RANDOM}};
  DMemory_1016 = _RAND_1054[31:0];
  _RAND_1055 = {1{`RANDOM}};
  DMemory_1017 = _RAND_1055[31:0];
  _RAND_1056 = {1{`RANDOM}};
  DMemory_1018 = _RAND_1056[31:0];
  _RAND_1057 = {1{`RANDOM}};
  DMemory_1019 = _RAND_1057[31:0];
  _RAND_1058 = {1{`RANDOM}};
  DMemory_1020 = _RAND_1058[31:0];
  _RAND_1059 = {1{`RANDOM}};
  DMemory_1021 = _RAND_1059[31:0];
  _RAND_1060 = {1{`RANDOM}};
  DMemory_1022 = _RAND_1060[31:0];
  _RAND_1061 = {1{`RANDOM}};
  DMemory_1023 = _RAND_1061[31:0];
  _RAND_1062 = {1{`RANDOM}};
  IMemory_0 = _RAND_1062[31:0];
  _RAND_1063 = {1{`RANDOM}};
  IMemory_1 = _RAND_1063[31:0];
  _RAND_1064 = {1{`RANDOM}};
  IMemory_2 = _RAND_1064[31:0];
  _RAND_1065 = {1{`RANDOM}};
  IMemory_3 = _RAND_1065[31:0];
  _RAND_1066 = {1{`RANDOM}};
  IMemory_4 = _RAND_1066[31:0];
  _RAND_1067 = {1{`RANDOM}};
  IMemory_5 = _RAND_1067[31:0];
  _RAND_1068 = {1{`RANDOM}};
  IMemory_6 = _RAND_1068[31:0];
  _RAND_1069 = {1{`RANDOM}};
  IMemory_7 = _RAND_1069[31:0];
  _RAND_1070 = {1{`RANDOM}};
  IFIDIR = _RAND_1070[31:0];
  _RAND_1071 = {1{`RANDOM}};
  IDEXIR = _RAND_1071[31:0];
  _RAND_1072 = {1{`RANDOM}};
  EXMEMIR = _RAND_1072[31:0];
  _RAND_1073 = {1{`RANDOM}};
  MEMWBIR = _RAND_1073[31:0];
  _RAND_1074 = {2{`RANDOM}};
  CurPC = _RAND_1074[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
