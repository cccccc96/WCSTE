module CAMLine(
  input         clock,
  input         io_we,
  input         io_wi,
  input  [63:0] io_key,
  input  [63:0] io_din,
  output        io_hit
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  write = io_we & io_wi; // @[cam.scala 58:18]
  reg [63:0] camCells; // @[cam.scala 59:21]
  assign io_hit = camCells == io_key; // @[cam.scala 65:23]
  always @(posedge clock) begin
    if (write) begin // @[cam.scala 61:14]
      camCells <= io_din; // @[cam.scala 62:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  camCells = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CAM_m_n(
  input         clock,
  input         reset,
  input         io_we,
  input  [63:0] io_key,
  input  [63:0] io_din,
  input  [63:0] io_waddr,
  output        io_hit
);
  wire  CAMLine_clock; // @[cam.scala 81:36]
  wire  CAMLine_io_we; // @[cam.scala 81:36]
  wire  CAMLine_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_io_din; // @[cam.scala 81:36]
  wire  CAMLine_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_1_clock; // @[cam.scala 81:36]
  wire  CAMLine_1_io_we; // @[cam.scala 81:36]
  wire  CAMLine_1_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_1_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_1_io_din; // @[cam.scala 81:36]
  wire  CAMLine_1_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_2_clock; // @[cam.scala 81:36]
  wire  CAMLine_2_io_we; // @[cam.scala 81:36]
  wire  CAMLine_2_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_2_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_2_io_din; // @[cam.scala 81:36]
  wire  CAMLine_2_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_3_clock; // @[cam.scala 81:36]
  wire  CAMLine_3_io_we; // @[cam.scala 81:36]
  wire  CAMLine_3_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_3_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_3_io_din; // @[cam.scala 81:36]
  wire  CAMLine_3_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_4_clock; // @[cam.scala 81:36]
  wire  CAMLine_4_io_we; // @[cam.scala 81:36]
  wire  CAMLine_4_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_4_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_4_io_din; // @[cam.scala 81:36]
  wire  CAMLine_4_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_5_clock; // @[cam.scala 81:36]
  wire  CAMLine_5_io_we; // @[cam.scala 81:36]
  wire  CAMLine_5_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_5_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_5_io_din; // @[cam.scala 81:36]
  wire  CAMLine_5_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_6_clock; // @[cam.scala 81:36]
  wire  CAMLine_6_io_we; // @[cam.scala 81:36]
  wire  CAMLine_6_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_6_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_6_io_din; // @[cam.scala 81:36]
  wire  CAMLine_6_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_7_clock; // @[cam.scala 81:36]
  wire  CAMLine_7_io_we; // @[cam.scala 81:36]
  wire  CAMLine_7_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_7_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_7_io_din; // @[cam.scala 81:36]
  wire  CAMLine_7_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_8_clock; // @[cam.scala 81:36]
  wire  CAMLine_8_io_we; // @[cam.scala 81:36]
  wire  CAMLine_8_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_8_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_8_io_din; // @[cam.scala 81:36]
  wire  CAMLine_8_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_9_clock; // @[cam.scala 81:36]
  wire  CAMLine_9_io_we; // @[cam.scala 81:36]
  wire  CAMLine_9_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_9_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_9_io_din; // @[cam.scala 81:36]
  wire  CAMLine_9_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_10_clock; // @[cam.scala 81:36]
  wire  CAMLine_10_io_we; // @[cam.scala 81:36]
  wire  CAMLine_10_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_10_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_10_io_din; // @[cam.scala 81:36]
  wire  CAMLine_10_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_11_clock; // @[cam.scala 81:36]
  wire  CAMLine_11_io_we; // @[cam.scala 81:36]
  wire  CAMLine_11_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_11_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_11_io_din; // @[cam.scala 81:36]
  wire  CAMLine_11_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_12_clock; // @[cam.scala 81:36]
  wire  CAMLine_12_io_we; // @[cam.scala 81:36]
  wire  CAMLine_12_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_12_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_12_io_din; // @[cam.scala 81:36]
  wire  CAMLine_12_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_13_clock; // @[cam.scala 81:36]
  wire  CAMLine_13_io_we; // @[cam.scala 81:36]
  wire  CAMLine_13_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_13_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_13_io_din; // @[cam.scala 81:36]
  wire  CAMLine_13_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_14_clock; // @[cam.scala 81:36]
  wire  CAMLine_14_io_we; // @[cam.scala 81:36]
  wire  CAMLine_14_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_14_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_14_io_din; // @[cam.scala 81:36]
  wire  CAMLine_14_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_15_clock; // @[cam.scala 81:36]
  wire  CAMLine_15_io_we; // @[cam.scala 81:36]
  wire  CAMLine_15_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_15_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_15_io_din; // @[cam.scala 81:36]
  wire  CAMLine_15_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_16_clock; // @[cam.scala 81:36]
  wire  CAMLine_16_io_we; // @[cam.scala 81:36]
  wire  CAMLine_16_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_16_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_16_io_din; // @[cam.scala 81:36]
  wire  CAMLine_16_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_17_clock; // @[cam.scala 81:36]
  wire  CAMLine_17_io_we; // @[cam.scala 81:36]
  wire  CAMLine_17_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_17_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_17_io_din; // @[cam.scala 81:36]
  wire  CAMLine_17_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_18_clock; // @[cam.scala 81:36]
  wire  CAMLine_18_io_we; // @[cam.scala 81:36]
  wire  CAMLine_18_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_18_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_18_io_din; // @[cam.scala 81:36]
  wire  CAMLine_18_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_19_clock; // @[cam.scala 81:36]
  wire  CAMLine_19_io_we; // @[cam.scala 81:36]
  wire  CAMLine_19_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_19_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_19_io_din; // @[cam.scala 81:36]
  wire  CAMLine_19_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_20_clock; // @[cam.scala 81:36]
  wire  CAMLine_20_io_we; // @[cam.scala 81:36]
  wire  CAMLine_20_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_20_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_20_io_din; // @[cam.scala 81:36]
  wire  CAMLine_20_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_21_clock; // @[cam.scala 81:36]
  wire  CAMLine_21_io_we; // @[cam.scala 81:36]
  wire  CAMLine_21_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_21_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_21_io_din; // @[cam.scala 81:36]
  wire  CAMLine_21_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_22_clock; // @[cam.scala 81:36]
  wire  CAMLine_22_io_we; // @[cam.scala 81:36]
  wire  CAMLine_22_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_22_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_22_io_din; // @[cam.scala 81:36]
  wire  CAMLine_22_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_23_clock; // @[cam.scala 81:36]
  wire  CAMLine_23_io_we; // @[cam.scala 81:36]
  wire  CAMLine_23_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_23_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_23_io_din; // @[cam.scala 81:36]
  wire  CAMLine_23_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_24_clock; // @[cam.scala 81:36]
  wire  CAMLine_24_io_we; // @[cam.scala 81:36]
  wire  CAMLine_24_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_24_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_24_io_din; // @[cam.scala 81:36]
  wire  CAMLine_24_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_25_clock; // @[cam.scala 81:36]
  wire  CAMLine_25_io_we; // @[cam.scala 81:36]
  wire  CAMLine_25_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_25_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_25_io_din; // @[cam.scala 81:36]
  wire  CAMLine_25_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_26_clock; // @[cam.scala 81:36]
  wire  CAMLine_26_io_we; // @[cam.scala 81:36]
  wire  CAMLine_26_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_26_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_26_io_din; // @[cam.scala 81:36]
  wire  CAMLine_26_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_27_clock; // @[cam.scala 81:36]
  wire  CAMLine_27_io_we; // @[cam.scala 81:36]
  wire  CAMLine_27_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_27_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_27_io_din; // @[cam.scala 81:36]
  wire  CAMLine_27_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_28_clock; // @[cam.scala 81:36]
  wire  CAMLine_28_io_we; // @[cam.scala 81:36]
  wire  CAMLine_28_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_28_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_28_io_din; // @[cam.scala 81:36]
  wire  CAMLine_28_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_29_clock; // @[cam.scala 81:36]
  wire  CAMLine_29_io_we; // @[cam.scala 81:36]
  wire  CAMLine_29_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_29_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_29_io_din; // @[cam.scala 81:36]
  wire  CAMLine_29_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_30_clock; // @[cam.scala 81:36]
  wire  CAMLine_30_io_we; // @[cam.scala 81:36]
  wire  CAMLine_30_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_30_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_30_io_din; // @[cam.scala 81:36]
  wire  CAMLine_30_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_31_clock; // @[cam.scala 81:36]
  wire  CAMLine_31_io_we; // @[cam.scala 81:36]
  wire  CAMLine_31_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_31_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_31_io_din; // @[cam.scala 81:36]
  wire  CAMLine_31_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_32_clock; // @[cam.scala 81:36]
  wire  CAMLine_32_io_we; // @[cam.scala 81:36]
  wire  CAMLine_32_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_32_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_32_io_din; // @[cam.scala 81:36]
  wire  CAMLine_32_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_33_clock; // @[cam.scala 81:36]
  wire  CAMLine_33_io_we; // @[cam.scala 81:36]
  wire  CAMLine_33_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_33_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_33_io_din; // @[cam.scala 81:36]
  wire  CAMLine_33_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_34_clock; // @[cam.scala 81:36]
  wire  CAMLine_34_io_we; // @[cam.scala 81:36]
  wire  CAMLine_34_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_34_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_34_io_din; // @[cam.scala 81:36]
  wire  CAMLine_34_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_35_clock; // @[cam.scala 81:36]
  wire  CAMLine_35_io_we; // @[cam.scala 81:36]
  wire  CAMLine_35_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_35_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_35_io_din; // @[cam.scala 81:36]
  wire  CAMLine_35_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_36_clock; // @[cam.scala 81:36]
  wire  CAMLine_36_io_we; // @[cam.scala 81:36]
  wire  CAMLine_36_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_36_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_36_io_din; // @[cam.scala 81:36]
  wire  CAMLine_36_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_37_clock; // @[cam.scala 81:36]
  wire  CAMLine_37_io_we; // @[cam.scala 81:36]
  wire  CAMLine_37_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_37_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_37_io_din; // @[cam.scala 81:36]
  wire  CAMLine_37_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_38_clock; // @[cam.scala 81:36]
  wire  CAMLine_38_io_we; // @[cam.scala 81:36]
  wire  CAMLine_38_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_38_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_38_io_din; // @[cam.scala 81:36]
  wire  CAMLine_38_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_39_clock; // @[cam.scala 81:36]
  wire  CAMLine_39_io_we; // @[cam.scala 81:36]
  wire  CAMLine_39_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_39_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_39_io_din; // @[cam.scala 81:36]
  wire  CAMLine_39_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_40_clock; // @[cam.scala 81:36]
  wire  CAMLine_40_io_we; // @[cam.scala 81:36]
  wire  CAMLine_40_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_40_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_40_io_din; // @[cam.scala 81:36]
  wire  CAMLine_40_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_41_clock; // @[cam.scala 81:36]
  wire  CAMLine_41_io_we; // @[cam.scala 81:36]
  wire  CAMLine_41_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_41_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_41_io_din; // @[cam.scala 81:36]
  wire  CAMLine_41_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_42_clock; // @[cam.scala 81:36]
  wire  CAMLine_42_io_we; // @[cam.scala 81:36]
  wire  CAMLine_42_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_42_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_42_io_din; // @[cam.scala 81:36]
  wire  CAMLine_42_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_43_clock; // @[cam.scala 81:36]
  wire  CAMLine_43_io_we; // @[cam.scala 81:36]
  wire  CAMLine_43_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_43_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_43_io_din; // @[cam.scala 81:36]
  wire  CAMLine_43_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_44_clock; // @[cam.scala 81:36]
  wire  CAMLine_44_io_we; // @[cam.scala 81:36]
  wire  CAMLine_44_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_44_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_44_io_din; // @[cam.scala 81:36]
  wire  CAMLine_44_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_45_clock; // @[cam.scala 81:36]
  wire  CAMLine_45_io_we; // @[cam.scala 81:36]
  wire  CAMLine_45_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_45_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_45_io_din; // @[cam.scala 81:36]
  wire  CAMLine_45_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_46_clock; // @[cam.scala 81:36]
  wire  CAMLine_46_io_we; // @[cam.scala 81:36]
  wire  CAMLine_46_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_46_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_46_io_din; // @[cam.scala 81:36]
  wire  CAMLine_46_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_47_clock; // @[cam.scala 81:36]
  wire  CAMLine_47_io_we; // @[cam.scala 81:36]
  wire  CAMLine_47_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_47_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_47_io_din; // @[cam.scala 81:36]
  wire  CAMLine_47_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_48_clock; // @[cam.scala 81:36]
  wire  CAMLine_48_io_we; // @[cam.scala 81:36]
  wire  CAMLine_48_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_48_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_48_io_din; // @[cam.scala 81:36]
  wire  CAMLine_48_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_49_clock; // @[cam.scala 81:36]
  wire  CAMLine_49_io_we; // @[cam.scala 81:36]
  wire  CAMLine_49_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_49_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_49_io_din; // @[cam.scala 81:36]
  wire  CAMLine_49_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_50_clock; // @[cam.scala 81:36]
  wire  CAMLine_50_io_we; // @[cam.scala 81:36]
  wire  CAMLine_50_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_50_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_50_io_din; // @[cam.scala 81:36]
  wire  CAMLine_50_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_51_clock; // @[cam.scala 81:36]
  wire  CAMLine_51_io_we; // @[cam.scala 81:36]
  wire  CAMLine_51_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_51_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_51_io_din; // @[cam.scala 81:36]
  wire  CAMLine_51_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_52_clock; // @[cam.scala 81:36]
  wire  CAMLine_52_io_we; // @[cam.scala 81:36]
  wire  CAMLine_52_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_52_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_52_io_din; // @[cam.scala 81:36]
  wire  CAMLine_52_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_53_clock; // @[cam.scala 81:36]
  wire  CAMLine_53_io_we; // @[cam.scala 81:36]
  wire  CAMLine_53_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_53_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_53_io_din; // @[cam.scala 81:36]
  wire  CAMLine_53_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_54_clock; // @[cam.scala 81:36]
  wire  CAMLine_54_io_we; // @[cam.scala 81:36]
  wire  CAMLine_54_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_54_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_54_io_din; // @[cam.scala 81:36]
  wire  CAMLine_54_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_55_clock; // @[cam.scala 81:36]
  wire  CAMLine_55_io_we; // @[cam.scala 81:36]
  wire  CAMLine_55_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_55_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_55_io_din; // @[cam.scala 81:36]
  wire  CAMLine_55_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_56_clock; // @[cam.scala 81:36]
  wire  CAMLine_56_io_we; // @[cam.scala 81:36]
  wire  CAMLine_56_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_56_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_56_io_din; // @[cam.scala 81:36]
  wire  CAMLine_56_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_57_clock; // @[cam.scala 81:36]
  wire  CAMLine_57_io_we; // @[cam.scala 81:36]
  wire  CAMLine_57_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_57_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_57_io_din; // @[cam.scala 81:36]
  wire  CAMLine_57_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_58_clock; // @[cam.scala 81:36]
  wire  CAMLine_58_io_we; // @[cam.scala 81:36]
  wire  CAMLine_58_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_58_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_58_io_din; // @[cam.scala 81:36]
  wire  CAMLine_58_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_59_clock; // @[cam.scala 81:36]
  wire  CAMLine_59_io_we; // @[cam.scala 81:36]
  wire  CAMLine_59_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_59_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_59_io_din; // @[cam.scala 81:36]
  wire  CAMLine_59_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_60_clock; // @[cam.scala 81:36]
  wire  CAMLine_60_io_we; // @[cam.scala 81:36]
  wire  CAMLine_60_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_60_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_60_io_din; // @[cam.scala 81:36]
  wire  CAMLine_60_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_61_clock; // @[cam.scala 81:36]
  wire  CAMLine_61_io_we; // @[cam.scala 81:36]
  wire  CAMLine_61_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_61_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_61_io_din; // @[cam.scala 81:36]
  wire  CAMLine_61_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_62_clock; // @[cam.scala 81:36]
  wire  CAMLine_62_io_we; // @[cam.scala 81:36]
  wire  CAMLine_62_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_62_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_62_io_din; // @[cam.scala 81:36]
  wire  CAMLine_62_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_63_clock; // @[cam.scala 81:36]
  wire  CAMLine_63_io_we; // @[cam.scala 81:36]
  wire  CAMLine_63_io_wi; // @[cam.scala 81:36]
  wire [63:0] CAMLine_63_io_key; // @[cam.scala 81:36]
  wire [63:0] CAMLine_63_io_din; // @[cam.scala 81:36]
  wire  CAMLine_63_io_hit; // @[cam.scala 81:36]
  wire  _io_hit_T_29 = CAMLine_io_hit | CAMLine_1_io_hit | CAMLine_2_io_hit | CAMLine_3_io_hit | CAMLine_4_io_hit |
    CAMLine_5_io_hit | CAMLine_6_io_hit | CAMLine_7_io_hit | CAMLine_8_io_hit | CAMLine_9_io_hit | CAMLine_10_io_hit |
    CAMLine_11_io_hit | CAMLine_12_io_hit | CAMLine_13_io_hit | CAMLine_14_io_hit | CAMLine_15_io_hit |
    CAMLine_16_io_hit | CAMLine_17_io_hit | CAMLine_18_io_hit | CAMLine_19_io_hit | CAMLine_20_io_hit |
    CAMLine_21_io_hit | CAMLine_22_io_hit | CAMLine_23_io_hit | CAMLine_24_io_hit | CAMLine_25_io_hit |
    CAMLine_26_io_hit | CAMLine_27_io_hit | CAMLine_28_io_hit | CAMLine_29_io_hit | CAMLine_30_io_hit; // @[cam.scala 93:27]
  wire  _io_hit_T_59 = _io_hit_T_29 | CAMLine_31_io_hit | CAMLine_32_io_hit | CAMLine_33_io_hit | CAMLine_34_io_hit |
    CAMLine_35_io_hit | CAMLine_36_io_hit | CAMLine_37_io_hit | CAMLine_38_io_hit | CAMLine_39_io_hit |
    CAMLine_40_io_hit | CAMLine_41_io_hit | CAMLine_42_io_hit | CAMLine_43_io_hit | CAMLine_44_io_hit |
    CAMLine_45_io_hit | CAMLine_46_io_hit | CAMLine_47_io_hit | CAMLine_48_io_hit | CAMLine_49_io_hit |
    CAMLine_50_io_hit | CAMLine_51_io_hit | CAMLine_52_io_hit | CAMLine_53_io_hit | CAMLine_54_io_hit |
    CAMLine_55_io_hit | CAMLine_56_io_hit | CAMLine_57_io_hit | CAMLine_58_io_hit | CAMLine_59_io_hit |
    CAMLine_60_io_hit; // @[cam.scala 93:27]
  CAMLine CAMLine ( // @[cam.scala 81:36]
    .clock(CAMLine_clock),
    .io_we(CAMLine_io_we),
    .io_wi(CAMLine_io_wi),
    .io_key(CAMLine_io_key),
    .io_din(CAMLine_io_din),
    .io_hit(CAMLine_io_hit)
  );
  CAMLine CAMLine_1 ( // @[cam.scala 81:36]
    .clock(CAMLine_1_clock),
    .io_we(CAMLine_1_io_we),
    .io_wi(CAMLine_1_io_wi),
    .io_key(CAMLine_1_io_key),
    .io_din(CAMLine_1_io_din),
    .io_hit(CAMLine_1_io_hit)
  );
  CAMLine CAMLine_2 ( // @[cam.scala 81:36]
    .clock(CAMLine_2_clock),
    .io_we(CAMLine_2_io_we),
    .io_wi(CAMLine_2_io_wi),
    .io_key(CAMLine_2_io_key),
    .io_din(CAMLine_2_io_din),
    .io_hit(CAMLine_2_io_hit)
  );
  CAMLine CAMLine_3 ( // @[cam.scala 81:36]
    .clock(CAMLine_3_clock),
    .io_we(CAMLine_3_io_we),
    .io_wi(CAMLine_3_io_wi),
    .io_key(CAMLine_3_io_key),
    .io_din(CAMLine_3_io_din),
    .io_hit(CAMLine_3_io_hit)
  );
  CAMLine CAMLine_4 ( // @[cam.scala 81:36]
    .clock(CAMLine_4_clock),
    .io_we(CAMLine_4_io_we),
    .io_wi(CAMLine_4_io_wi),
    .io_key(CAMLine_4_io_key),
    .io_din(CAMLine_4_io_din),
    .io_hit(CAMLine_4_io_hit)
  );
  CAMLine CAMLine_5 ( // @[cam.scala 81:36]
    .clock(CAMLine_5_clock),
    .io_we(CAMLine_5_io_we),
    .io_wi(CAMLine_5_io_wi),
    .io_key(CAMLine_5_io_key),
    .io_din(CAMLine_5_io_din),
    .io_hit(CAMLine_5_io_hit)
  );
  CAMLine CAMLine_6 ( // @[cam.scala 81:36]
    .clock(CAMLine_6_clock),
    .io_we(CAMLine_6_io_we),
    .io_wi(CAMLine_6_io_wi),
    .io_key(CAMLine_6_io_key),
    .io_din(CAMLine_6_io_din),
    .io_hit(CAMLine_6_io_hit)
  );
  CAMLine CAMLine_7 ( // @[cam.scala 81:36]
    .clock(CAMLine_7_clock),
    .io_we(CAMLine_7_io_we),
    .io_wi(CAMLine_7_io_wi),
    .io_key(CAMLine_7_io_key),
    .io_din(CAMLine_7_io_din),
    .io_hit(CAMLine_7_io_hit)
  );
  CAMLine CAMLine_8 ( // @[cam.scala 81:36]
    .clock(CAMLine_8_clock),
    .io_we(CAMLine_8_io_we),
    .io_wi(CAMLine_8_io_wi),
    .io_key(CAMLine_8_io_key),
    .io_din(CAMLine_8_io_din),
    .io_hit(CAMLine_8_io_hit)
  );
  CAMLine CAMLine_9 ( // @[cam.scala 81:36]
    .clock(CAMLine_9_clock),
    .io_we(CAMLine_9_io_we),
    .io_wi(CAMLine_9_io_wi),
    .io_key(CAMLine_9_io_key),
    .io_din(CAMLine_9_io_din),
    .io_hit(CAMLine_9_io_hit)
  );
  CAMLine CAMLine_10 ( // @[cam.scala 81:36]
    .clock(CAMLine_10_clock),
    .io_we(CAMLine_10_io_we),
    .io_wi(CAMLine_10_io_wi),
    .io_key(CAMLine_10_io_key),
    .io_din(CAMLine_10_io_din),
    .io_hit(CAMLine_10_io_hit)
  );
  CAMLine CAMLine_11 ( // @[cam.scala 81:36]
    .clock(CAMLine_11_clock),
    .io_we(CAMLine_11_io_we),
    .io_wi(CAMLine_11_io_wi),
    .io_key(CAMLine_11_io_key),
    .io_din(CAMLine_11_io_din),
    .io_hit(CAMLine_11_io_hit)
  );
  CAMLine CAMLine_12 ( // @[cam.scala 81:36]
    .clock(CAMLine_12_clock),
    .io_we(CAMLine_12_io_we),
    .io_wi(CAMLine_12_io_wi),
    .io_key(CAMLine_12_io_key),
    .io_din(CAMLine_12_io_din),
    .io_hit(CAMLine_12_io_hit)
  );
  CAMLine CAMLine_13 ( // @[cam.scala 81:36]
    .clock(CAMLine_13_clock),
    .io_we(CAMLine_13_io_we),
    .io_wi(CAMLine_13_io_wi),
    .io_key(CAMLine_13_io_key),
    .io_din(CAMLine_13_io_din),
    .io_hit(CAMLine_13_io_hit)
  );
  CAMLine CAMLine_14 ( // @[cam.scala 81:36]
    .clock(CAMLine_14_clock),
    .io_we(CAMLine_14_io_we),
    .io_wi(CAMLine_14_io_wi),
    .io_key(CAMLine_14_io_key),
    .io_din(CAMLine_14_io_din),
    .io_hit(CAMLine_14_io_hit)
  );
  CAMLine CAMLine_15 ( // @[cam.scala 81:36]
    .clock(CAMLine_15_clock),
    .io_we(CAMLine_15_io_we),
    .io_wi(CAMLine_15_io_wi),
    .io_key(CAMLine_15_io_key),
    .io_din(CAMLine_15_io_din),
    .io_hit(CAMLine_15_io_hit)
  );
  CAMLine CAMLine_16 ( // @[cam.scala 81:36]
    .clock(CAMLine_16_clock),
    .io_we(CAMLine_16_io_we),
    .io_wi(CAMLine_16_io_wi),
    .io_key(CAMLine_16_io_key),
    .io_din(CAMLine_16_io_din),
    .io_hit(CAMLine_16_io_hit)
  );
  CAMLine CAMLine_17 ( // @[cam.scala 81:36]
    .clock(CAMLine_17_clock),
    .io_we(CAMLine_17_io_we),
    .io_wi(CAMLine_17_io_wi),
    .io_key(CAMLine_17_io_key),
    .io_din(CAMLine_17_io_din),
    .io_hit(CAMLine_17_io_hit)
  );
  CAMLine CAMLine_18 ( // @[cam.scala 81:36]
    .clock(CAMLine_18_clock),
    .io_we(CAMLine_18_io_we),
    .io_wi(CAMLine_18_io_wi),
    .io_key(CAMLine_18_io_key),
    .io_din(CAMLine_18_io_din),
    .io_hit(CAMLine_18_io_hit)
  );
  CAMLine CAMLine_19 ( // @[cam.scala 81:36]
    .clock(CAMLine_19_clock),
    .io_we(CAMLine_19_io_we),
    .io_wi(CAMLine_19_io_wi),
    .io_key(CAMLine_19_io_key),
    .io_din(CAMLine_19_io_din),
    .io_hit(CAMLine_19_io_hit)
  );
  CAMLine CAMLine_20 ( // @[cam.scala 81:36]
    .clock(CAMLine_20_clock),
    .io_we(CAMLine_20_io_we),
    .io_wi(CAMLine_20_io_wi),
    .io_key(CAMLine_20_io_key),
    .io_din(CAMLine_20_io_din),
    .io_hit(CAMLine_20_io_hit)
  );
  CAMLine CAMLine_21 ( // @[cam.scala 81:36]
    .clock(CAMLine_21_clock),
    .io_we(CAMLine_21_io_we),
    .io_wi(CAMLine_21_io_wi),
    .io_key(CAMLine_21_io_key),
    .io_din(CAMLine_21_io_din),
    .io_hit(CAMLine_21_io_hit)
  );
  CAMLine CAMLine_22 ( // @[cam.scala 81:36]
    .clock(CAMLine_22_clock),
    .io_we(CAMLine_22_io_we),
    .io_wi(CAMLine_22_io_wi),
    .io_key(CAMLine_22_io_key),
    .io_din(CAMLine_22_io_din),
    .io_hit(CAMLine_22_io_hit)
  );
  CAMLine CAMLine_23 ( // @[cam.scala 81:36]
    .clock(CAMLine_23_clock),
    .io_we(CAMLine_23_io_we),
    .io_wi(CAMLine_23_io_wi),
    .io_key(CAMLine_23_io_key),
    .io_din(CAMLine_23_io_din),
    .io_hit(CAMLine_23_io_hit)
  );
  CAMLine CAMLine_24 ( // @[cam.scala 81:36]
    .clock(CAMLine_24_clock),
    .io_we(CAMLine_24_io_we),
    .io_wi(CAMLine_24_io_wi),
    .io_key(CAMLine_24_io_key),
    .io_din(CAMLine_24_io_din),
    .io_hit(CAMLine_24_io_hit)
  );
  CAMLine CAMLine_25 ( // @[cam.scala 81:36]
    .clock(CAMLine_25_clock),
    .io_we(CAMLine_25_io_we),
    .io_wi(CAMLine_25_io_wi),
    .io_key(CAMLine_25_io_key),
    .io_din(CAMLine_25_io_din),
    .io_hit(CAMLine_25_io_hit)
  );
  CAMLine CAMLine_26 ( // @[cam.scala 81:36]
    .clock(CAMLine_26_clock),
    .io_we(CAMLine_26_io_we),
    .io_wi(CAMLine_26_io_wi),
    .io_key(CAMLine_26_io_key),
    .io_din(CAMLine_26_io_din),
    .io_hit(CAMLine_26_io_hit)
  );
  CAMLine CAMLine_27 ( // @[cam.scala 81:36]
    .clock(CAMLine_27_clock),
    .io_we(CAMLine_27_io_we),
    .io_wi(CAMLine_27_io_wi),
    .io_key(CAMLine_27_io_key),
    .io_din(CAMLine_27_io_din),
    .io_hit(CAMLine_27_io_hit)
  );
  CAMLine CAMLine_28 ( // @[cam.scala 81:36]
    .clock(CAMLine_28_clock),
    .io_we(CAMLine_28_io_we),
    .io_wi(CAMLine_28_io_wi),
    .io_key(CAMLine_28_io_key),
    .io_din(CAMLine_28_io_din),
    .io_hit(CAMLine_28_io_hit)
  );
  CAMLine CAMLine_29 ( // @[cam.scala 81:36]
    .clock(CAMLine_29_clock),
    .io_we(CAMLine_29_io_we),
    .io_wi(CAMLine_29_io_wi),
    .io_key(CAMLine_29_io_key),
    .io_din(CAMLine_29_io_din),
    .io_hit(CAMLine_29_io_hit)
  );
  CAMLine CAMLine_30 ( // @[cam.scala 81:36]
    .clock(CAMLine_30_clock),
    .io_we(CAMLine_30_io_we),
    .io_wi(CAMLine_30_io_wi),
    .io_key(CAMLine_30_io_key),
    .io_din(CAMLine_30_io_din),
    .io_hit(CAMLine_30_io_hit)
  );
  CAMLine CAMLine_31 ( // @[cam.scala 81:36]
    .clock(CAMLine_31_clock),
    .io_we(CAMLine_31_io_we),
    .io_wi(CAMLine_31_io_wi),
    .io_key(CAMLine_31_io_key),
    .io_din(CAMLine_31_io_din),
    .io_hit(CAMLine_31_io_hit)
  );
  CAMLine CAMLine_32 ( // @[cam.scala 81:36]
    .clock(CAMLine_32_clock),
    .io_we(CAMLine_32_io_we),
    .io_wi(CAMLine_32_io_wi),
    .io_key(CAMLine_32_io_key),
    .io_din(CAMLine_32_io_din),
    .io_hit(CAMLine_32_io_hit)
  );
  CAMLine CAMLine_33 ( // @[cam.scala 81:36]
    .clock(CAMLine_33_clock),
    .io_we(CAMLine_33_io_we),
    .io_wi(CAMLine_33_io_wi),
    .io_key(CAMLine_33_io_key),
    .io_din(CAMLine_33_io_din),
    .io_hit(CAMLine_33_io_hit)
  );
  CAMLine CAMLine_34 ( // @[cam.scala 81:36]
    .clock(CAMLine_34_clock),
    .io_we(CAMLine_34_io_we),
    .io_wi(CAMLine_34_io_wi),
    .io_key(CAMLine_34_io_key),
    .io_din(CAMLine_34_io_din),
    .io_hit(CAMLine_34_io_hit)
  );
  CAMLine CAMLine_35 ( // @[cam.scala 81:36]
    .clock(CAMLine_35_clock),
    .io_we(CAMLine_35_io_we),
    .io_wi(CAMLine_35_io_wi),
    .io_key(CAMLine_35_io_key),
    .io_din(CAMLine_35_io_din),
    .io_hit(CAMLine_35_io_hit)
  );
  CAMLine CAMLine_36 ( // @[cam.scala 81:36]
    .clock(CAMLine_36_clock),
    .io_we(CAMLine_36_io_we),
    .io_wi(CAMLine_36_io_wi),
    .io_key(CAMLine_36_io_key),
    .io_din(CAMLine_36_io_din),
    .io_hit(CAMLine_36_io_hit)
  );
  CAMLine CAMLine_37 ( // @[cam.scala 81:36]
    .clock(CAMLine_37_clock),
    .io_we(CAMLine_37_io_we),
    .io_wi(CAMLine_37_io_wi),
    .io_key(CAMLine_37_io_key),
    .io_din(CAMLine_37_io_din),
    .io_hit(CAMLine_37_io_hit)
  );
  CAMLine CAMLine_38 ( // @[cam.scala 81:36]
    .clock(CAMLine_38_clock),
    .io_we(CAMLine_38_io_we),
    .io_wi(CAMLine_38_io_wi),
    .io_key(CAMLine_38_io_key),
    .io_din(CAMLine_38_io_din),
    .io_hit(CAMLine_38_io_hit)
  );
  CAMLine CAMLine_39 ( // @[cam.scala 81:36]
    .clock(CAMLine_39_clock),
    .io_we(CAMLine_39_io_we),
    .io_wi(CAMLine_39_io_wi),
    .io_key(CAMLine_39_io_key),
    .io_din(CAMLine_39_io_din),
    .io_hit(CAMLine_39_io_hit)
  );
  CAMLine CAMLine_40 ( // @[cam.scala 81:36]
    .clock(CAMLine_40_clock),
    .io_we(CAMLine_40_io_we),
    .io_wi(CAMLine_40_io_wi),
    .io_key(CAMLine_40_io_key),
    .io_din(CAMLine_40_io_din),
    .io_hit(CAMLine_40_io_hit)
  );
  CAMLine CAMLine_41 ( // @[cam.scala 81:36]
    .clock(CAMLine_41_clock),
    .io_we(CAMLine_41_io_we),
    .io_wi(CAMLine_41_io_wi),
    .io_key(CAMLine_41_io_key),
    .io_din(CAMLine_41_io_din),
    .io_hit(CAMLine_41_io_hit)
  );
  CAMLine CAMLine_42 ( // @[cam.scala 81:36]
    .clock(CAMLine_42_clock),
    .io_we(CAMLine_42_io_we),
    .io_wi(CAMLine_42_io_wi),
    .io_key(CAMLine_42_io_key),
    .io_din(CAMLine_42_io_din),
    .io_hit(CAMLine_42_io_hit)
  );
  CAMLine CAMLine_43 ( // @[cam.scala 81:36]
    .clock(CAMLine_43_clock),
    .io_we(CAMLine_43_io_we),
    .io_wi(CAMLine_43_io_wi),
    .io_key(CAMLine_43_io_key),
    .io_din(CAMLine_43_io_din),
    .io_hit(CAMLine_43_io_hit)
  );
  CAMLine CAMLine_44 ( // @[cam.scala 81:36]
    .clock(CAMLine_44_clock),
    .io_we(CAMLine_44_io_we),
    .io_wi(CAMLine_44_io_wi),
    .io_key(CAMLine_44_io_key),
    .io_din(CAMLine_44_io_din),
    .io_hit(CAMLine_44_io_hit)
  );
  CAMLine CAMLine_45 ( // @[cam.scala 81:36]
    .clock(CAMLine_45_clock),
    .io_we(CAMLine_45_io_we),
    .io_wi(CAMLine_45_io_wi),
    .io_key(CAMLine_45_io_key),
    .io_din(CAMLine_45_io_din),
    .io_hit(CAMLine_45_io_hit)
  );
  CAMLine CAMLine_46 ( // @[cam.scala 81:36]
    .clock(CAMLine_46_clock),
    .io_we(CAMLine_46_io_we),
    .io_wi(CAMLine_46_io_wi),
    .io_key(CAMLine_46_io_key),
    .io_din(CAMLine_46_io_din),
    .io_hit(CAMLine_46_io_hit)
  );
  CAMLine CAMLine_47 ( // @[cam.scala 81:36]
    .clock(CAMLine_47_clock),
    .io_we(CAMLine_47_io_we),
    .io_wi(CAMLine_47_io_wi),
    .io_key(CAMLine_47_io_key),
    .io_din(CAMLine_47_io_din),
    .io_hit(CAMLine_47_io_hit)
  );
  CAMLine CAMLine_48 ( // @[cam.scala 81:36]
    .clock(CAMLine_48_clock),
    .io_we(CAMLine_48_io_we),
    .io_wi(CAMLine_48_io_wi),
    .io_key(CAMLine_48_io_key),
    .io_din(CAMLine_48_io_din),
    .io_hit(CAMLine_48_io_hit)
  );
  CAMLine CAMLine_49 ( // @[cam.scala 81:36]
    .clock(CAMLine_49_clock),
    .io_we(CAMLine_49_io_we),
    .io_wi(CAMLine_49_io_wi),
    .io_key(CAMLine_49_io_key),
    .io_din(CAMLine_49_io_din),
    .io_hit(CAMLine_49_io_hit)
  );
  CAMLine CAMLine_50 ( // @[cam.scala 81:36]
    .clock(CAMLine_50_clock),
    .io_we(CAMLine_50_io_we),
    .io_wi(CAMLine_50_io_wi),
    .io_key(CAMLine_50_io_key),
    .io_din(CAMLine_50_io_din),
    .io_hit(CAMLine_50_io_hit)
  );
  CAMLine CAMLine_51 ( // @[cam.scala 81:36]
    .clock(CAMLine_51_clock),
    .io_we(CAMLine_51_io_we),
    .io_wi(CAMLine_51_io_wi),
    .io_key(CAMLine_51_io_key),
    .io_din(CAMLine_51_io_din),
    .io_hit(CAMLine_51_io_hit)
  );
  CAMLine CAMLine_52 ( // @[cam.scala 81:36]
    .clock(CAMLine_52_clock),
    .io_we(CAMLine_52_io_we),
    .io_wi(CAMLine_52_io_wi),
    .io_key(CAMLine_52_io_key),
    .io_din(CAMLine_52_io_din),
    .io_hit(CAMLine_52_io_hit)
  );
  CAMLine CAMLine_53 ( // @[cam.scala 81:36]
    .clock(CAMLine_53_clock),
    .io_we(CAMLine_53_io_we),
    .io_wi(CAMLine_53_io_wi),
    .io_key(CAMLine_53_io_key),
    .io_din(CAMLine_53_io_din),
    .io_hit(CAMLine_53_io_hit)
  );
  CAMLine CAMLine_54 ( // @[cam.scala 81:36]
    .clock(CAMLine_54_clock),
    .io_we(CAMLine_54_io_we),
    .io_wi(CAMLine_54_io_wi),
    .io_key(CAMLine_54_io_key),
    .io_din(CAMLine_54_io_din),
    .io_hit(CAMLine_54_io_hit)
  );
  CAMLine CAMLine_55 ( // @[cam.scala 81:36]
    .clock(CAMLine_55_clock),
    .io_we(CAMLine_55_io_we),
    .io_wi(CAMLine_55_io_wi),
    .io_key(CAMLine_55_io_key),
    .io_din(CAMLine_55_io_din),
    .io_hit(CAMLine_55_io_hit)
  );
  CAMLine CAMLine_56 ( // @[cam.scala 81:36]
    .clock(CAMLine_56_clock),
    .io_we(CAMLine_56_io_we),
    .io_wi(CAMLine_56_io_wi),
    .io_key(CAMLine_56_io_key),
    .io_din(CAMLine_56_io_din),
    .io_hit(CAMLine_56_io_hit)
  );
  CAMLine CAMLine_57 ( // @[cam.scala 81:36]
    .clock(CAMLine_57_clock),
    .io_we(CAMLine_57_io_we),
    .io_wi(CAMLine_57_io_wi),
    .io_key(CAMLine_57_io_key),
    .io_din(CAMLine_57_io_din),
    .io_hit(CAMLine_57_io_hit)
  );
  CAMLine CAMLine_58 ( // @[cam.scala 81:36]
    .clock(CAMLine_58_clock),
    .io_we(CAMLine_58_io_we),
    .io_wi(CAMLine_58_io_wi),
    .io_key(CAMLine_58_io_key),
    .io_din(CAMLine_58_io_din),
    .io_hit(CAMLine_58_io_hit)
  );
  CAMLine CAMLine_59 ( // @[cam.scala 81:36]
    .clock(CAMLine_59_clock),
    .io_we(CAMLine_59_io_we),
    .io_wi(CAMLine_59_io_wi),
    .io_key(CAMLine_59_io_key),
    .io_din(CAMLine_59_io_din),
    .io_hit(CAMLine_59_io_hit)
  );
  CAMLine CAMLine_60 ( // @[cam.scala 81:36]
    .clock(CAMLine_60_clock),
    .io_we(CAMLine_60_io_we),
    .io_wi(CAMLine_60_io_wi),
    .io_key(CAMLine_60_io_key),
    .io_din(CAMLine_60_io_din),
    .io_hit(CAMLine_60_io_hit)
  );
  CAMLine CAMLine_61 ( // @[cam.scala 81:36]
    .clock(CAMLine_61_clock),
    .io_we(CAMLine_61_io_we),
    .io_wi(CAMLine_61_io_wi),
    .io_key(CAMLine_61_io_key),
    .io_din(CAMLine_61_io_din),
    .io_hit(CAMLine_61_io_hit)
  );
  CAMLine CAMLine_62 ( // @[cam.scala 81:36]
    .clock(CAMLine_62_clock),
    .io_we(CAMLine_62_io_we),
    .io_wi(CAMLine_62_io_wi),
    .io_key(CAMLine_62_io_key),
    .io_din(CAMLine_62_io_din),
    .io_hit(CAMLine_62_io_hit)
  );
  CAMLine CAMLine_63 ( // @[cam.scala 81:36]
    .clock(CAMLine_63_clock),
    .io_we(CAMLine_63_io_we),
    .io_wi(CAMLine_63_io_wi),
    .io_key(CAMLine_63_io_key),
    .io_din(CAMLine_63_io_din),
    .io_hit(CAMLine_63_io_hit)
  );
  assign io_hit = _io_hit_T_59 | CAMLine_61_io_hit | CAMLine_62_io_hit | CAMLine_63_io_hit; // @[cam.scala 93:27]
  assign CAMLine_clock = clock;
  assign CAMLine_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_io_wi = io_waddr[0]; // @[cam.scala 86:31]
  assign CAMLine_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_1_clock = clock;
  assign CAMLine_1_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_1_io_wi = io_waddr[1]; // @[cam.scala 86:31]
  assign CAMLine_1_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_1_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_2_clock = clock;
  assign CAMLine_2_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_2_io_wi = io_waddr[2]; // @[cam.scala 86:31]
  assign CAMLine_2_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_2_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_3_clock = clock;
  assign CAMLine_3_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_3_io_wi = io_waddr[3]; // @[cam.scala 86:31]
  assign CAMLine_3_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_3_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_4_clock = clock;
  assign CAMLine_4_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_4_io_wi = io_waddr[4]; // @[cam.scala 86:31]
  assign CAMLine_4_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_4_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_5_clock = clock;
  assign CAMLine_5_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_5_io_wi = io_waddr[5]; // @[cam.scala 86:31]
  assign CAMLine_5_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_5_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_6_clock = clock;
  assign CAMLine_6_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_6_io_wi = io_waddr[6]; // @[cam.scala 86:31]
  assign CAMLine_6_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_6_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_7_clock = clock;
  assign CAMLine_7_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_7_io_wi = io_waddr[7]; // @[cam.scala 86:31]
  assign CAMLine_7_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_7_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_8_clock = clock;
  assign CAMLine_8_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_8_io_wi = io_waddr[8]; // @[cam.scala 86:31]
  assign CAMLine_8_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_8_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_9_clock = clock;
  assign CAMLine_9_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_9_io_wi = io_waddr[9]; // @[cam.scala 86:31]
  assign CAMLine_9_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_9_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_10_clock = clock;
  assign CAMLine_10_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_10_io_wi = io_waddr[10]; // @[cam.scala 86:31]
  assign CAMLine_10_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_10_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_11_clock = clock;
  assign CAMLine_11_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_11_io_wi = io_waddr[11]; // @[cam.scala 86:31]
  assign CAMLine_11_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_11_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_12_clock = clock;
  assign CAMLine_12_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_12_io_wi = io_waddr[12]; // @[cam.scala 86:31]
  assign CAMLine_12_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_12_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_13_clock = clock;
  assign CAMLine_13_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_13_io_wi = io_waddr[13]; // @[cam.scala 86:31]
  assign CAMLine_13_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_13_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_14_clock = clock;
  assign CAMLine_14_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_14_io_wi = io_waddr[14]; // @[cam.scala 86:31]
  assign CAMLine_14_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_14_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_15_clock = clock;
  assign CAMLine_15_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_15_io_wi = io_waddr[15]; // @[cam.scala 86:31]
  assign CAMLine_15_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_15_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_16_clock = clock;
  assign CAMLine_16_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_16_io_wi = io_waddr[16]; // @[cam.scala 86:31]
  assign CAMLine_16_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_16_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_17_clock = clock;
  assign CAMLine_17_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_17_io_wi = io_waddr[17]; // @[cam.scala 86:31]
  assign CAMLine_17_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_17_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_18_clock = clock;
  assign CAMLine_18_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_18_io_wi = io_waddr[18]; // @[cam.scala 86:31]
  assign CAMLine_18_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_18_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_19_clock = clock;
  assign CAMLine_19_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_19_io_wi = io_waddr[19]; // @[cam.scala 86:31]
  assign CAMLine_19_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_19_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_20_clock = clock;
  assign CAMLine_20_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_20_io_wi = io_waddr[20]; // @[cam.scala 86:31]
  assign CAMLine_20_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_20_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_21_clock = clock;
  assign CAMLine_21_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_21_io_wi = io_waddr[21]; // @[cam.scala 86:31]
  assign CAMLine_21_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_21_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_22_clock = clock;
  assign CAMLine_22_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_22_io_wi = io_waddr[22]; // @[cam.scala 86:31]
  assign CAMLine_22_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_22_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_23_clock = clock;
  assign CAMLine_23_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_23_io_wi = io_waddr[23]; // @[cam.scala 86:31]
  assign CAMLine_23_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_23_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_24_clock = clock;
  assign CAMLine_24_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_24_io_wi = io_waddr[24]; // @[cam.scala 86:31]
  assign CAMLine_24_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_24_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_25_clock = clock;
  assign CAMLine_25_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_25_io_wi = io_waddr[25]; // @[cam.scala 86:31]
  assign CAMLine_25_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_25_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_26_clock = clock;
  assign CAMLine_26_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_26_io_wi = io_waddr[26]; // @[cam.scala 86:31]
  assign CAMLine_26_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_26_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_27_clock = clock;
  assign CAMLine_27_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_27_io_wi = io_waddr[27]; // @[cam.scala 86:31]
  assign CAMLine_27_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_27_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_28_clock = clock;
  assign CAMLine_28_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_28_io_wi = io_waddr[28]; // @[cam.scala 86:31]
  assign CAMLine_28_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_28_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_29_clock = clock;
  assign CAMLine_29_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_29_io_wi = io_waddr[29]; // @[cam.scala 86:31]
  assign CAMLine_29_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_29_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_30_clock = clock;
  assign CAMLine_30_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_30_io_wi = io_waddr[30]; // @[cam.scala 86:31]
  assign CAMLine_30_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_30_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_31_clock = clock;
  assign CAMLine_31_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_31_io_wi = io_waddr[31]; // @[cam.scala 86:31]
  assign CAMLine_31_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_31_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_32_clock = clock;
  assign CAMLine_32_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_32_io_wi = io_waddr[32]; // @[cam.scala 86:31]
  assign CAMLine_32_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_32_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_33_clock = clock;
  assign CAMLine_33_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_33_io_wi = io_waddr[33]; // @[cam.scala 86:31]
  assign CAMLine_33_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_33_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_34_clock = clock;
  assign CAMLine_34_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_34_io_wi = io_waddr[34]; // @[cam.scala 86:31]
  assign CAMLine_34_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_34_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_35_clock = clock;
  assign CAMLine_35_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_35_io_wi = io_waddr[35]; // @[cam.scala 86:31]
  assign CAMLine_35_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_35_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_36_clock = clock;
  assign CAMLine_36_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_36_io_wi = io_waddr[36]; // @[cam.scala 86:31]
  assign CAMLine_36_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_36_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_37_clock = clock;
  assign CAMLine_37_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_37_io_wi = io_waddr[37]; // @[cam.scala 86:31]
  assign CAMLine_37_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_37_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_38_clock = clock;
  assign CAMLine_38_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_38_io_wi = io_waddr[38]; // @[cam.scala 86:31]
  assign CAMLine_38_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_38_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_39_clock = clock;
  assign CAMLine_39_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_39_io_wi = io_waddr[39]; // @[cam.scala 86:31]
  assign CAMLine_39_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_39_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_40_clock = clock;
  assign CAMLine_40_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_40_io_wi = io_waddr[40]; // @[cam.scala 86:31]
  assign CAMLine_40_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_40_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_41_clock = clock;
  assign CAMLine_41_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_41_io_wi = io_waddr[41]; // @[cam.scala 86:31]
  assign CAMLine_41_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_41_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_42_clock = clock;
  assign CAMLine_42_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_42_io_wi = io_waddr[42]; // @[cam.scala 86:31]
  assign CAMLine_42_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_42_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_43_clock = clock;
  assign CAMLine_43_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_43_io_wi = io_waddr[43]; // @[cam.scala 86:31]
  assign CAMLine_43_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_43_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_44_clock = clock;
  assign CAMLine_44_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_44_io_wi = io_waddr[44]; // @[cam.scala 86:31]
  assign CAMLine_44_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_44_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_45_clock = clock;
  assign CAMLine_45_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_45_io_wi = io_waddr[45]; // @[cam.scala 86:31]
  assign CAMLine_45_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_45_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_46_clock = clock;
  assign CAMLine_46_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_46_io_wi = io_waddr[46]; // @[cam.scala 86:31]
  assign CAMLine_46_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_46_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_47_clock = clock;
  assign CAMLine_47_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_47_io_wi = io_waddr[47]; // @[cam.scala 86:31]
  assign CAMLine_47_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_47_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_48_clock = clock;
  assign CAMLine_48_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_48_io_wi = io_waddr[48]; // @[cam.scala 86:31]
  assign CAMLine_48_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_48_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_49_clock = clock;
  assign CAMLine_49_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_49_io_wi = io_waddr[49]; // @[cam.scala 86:31]
  assign CAMLine_49_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_49_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_50_clock = clock;
  assign CAMLine_50_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_50_io_wi = io_waddr[50]; // @[cam.scala 86:31]
  assign CAMLine_50_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_50_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_51_clock = clock;
  assign CAMLine_51_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_51_io_wi = io_waddr[51]; // @[cam.scala 86:31]
  assign CAMLine_51_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_51_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_52_clock = clock;
  assign CAMLine_52_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_52_io_wi = io_waddr[52]; // @[cam.scala 86:31]
  assign CAMLine_52_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_52_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_53_clock = clock;
  assign CAMLine_53_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_53_io_wi = io_waddr[53]; // @[cam.scala 86:31]
  assign CAMLine_53_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_53_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_54_clock = clock;
  assign CAMLine_54_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_54_io_wi = io_waddr[54]; // @[cam.scala 86:31]
  assign CAMLine_54_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_54_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_55_clock = clock;
  assign CAMLine_55_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_55_io_wi = io_waddr[55]; // @[cam.scala 86:31]
  assign CAMLine_55_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_55_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_56_clock = clock;
  assign CAMLine_56_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_56_io_wi = io_waddr[56]; // @[cam.scala 86:31]
  assign CAMLine_56_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_56_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_57_clock = clock;
  assign CAMLine_57_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_57_io_wi = io_waddr[57]; // @[cam.scala 86:31]
  assign CAMLine_57_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_57_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_58_clock = clock;
  assign CAMLine_58_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_58_io_wi = io_waddr[58]; // @[cam.scala 86:31]
  assign CAMLine_58_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_58_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_59_clock = clock;
  assign CAMLine_59_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_59_io_wi = io_waddr[59]; // @[cam.scala 86:31]
  assign CAMLine_59_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_59_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_60_clock = clock;
  assign CAMLine_60_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_60_io_wi = io_waddr[60]; // @[cam.scala 86:31]
  assign CAMLine_60_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_60_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_61_clock = clock;
  assign CAMLine_61_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_61_io_wi = io_waddr[61]; // @[cam.scala 86:31]
  assign CAMLine_61_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_61_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_62_clock = clock;
  assign CAMLine_62_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_62_io_wi = io_waddr[62]; // @[cam.scala 86:31]
  assign CAMLine_62_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_62_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_63_clock = clock;
  assign CAMLine_63_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_63_io_wi = io_waddr[63]; // @[cam.scala 86:31]
  assign CAMLine_63_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_63_io_din = io_din; // @[cam.scala 88:21]
endmodule
