module RISCVCPUv2(
  input         clock,
  input         reset,
  input         io_rvfi_rst,
  input  [31:0] io_rvfi_insn_in_0,
  input  [31:0] io_rvfi_insn_in_1,
  output [63:0] io_rvfi_regs_0,
  output [63:0] io_rvfi_regs_1,
  output [63:0] io_rvfi_regs_2,
  output [63:0] io_rvfi_regs_3,
  output [63:0] io_rvfi_regs_4,
  output [63:0] io_rvfi_regs_5,
  output [63:0] io_rvfi_regs_6,
  output [63:0] io_rvfi_regs_7,
  output [63:0] io_rvfi_regs_8,
  output [63:0] io_rvfi_regs_9,
  output [63:0] io_rvfi_regs_10,
  output [63:0] io_rvfi_regs_11,
  output [63:0] io_rvfi_regs_12,
  output [63:0] io_rvfi_regs_13,
  output [63:0] io_rvfi_regs_14,
  output [63:0] io_rvfi_regs_15,
  output [63:0] io_rvfi_regs_16,
  output [63:0] io_rvfi_regs_17,
  output [63:0] io_rvfi_regs_18,
  output [63:0] io_rvfi_regs_19,
  output [63:0] io_rvfi_regs_20,
  output [63:0] io_rvfi_regs_21,
  output [63:0] io_rvfi_regs_22,
  output [63:0] io_rvfi_regs_23,
  output [63:0] io_rvfi_regs_24,
  output [63:0] io_rvfi_regs_25,
  output [63:0] io_rvfi_regs_26,
  output [63:0] io_rvfi_regs_27,
  output [63:0] io_rvfi_regs_28,
  output [63:0] io_rvfi_regs_29,
  output [63:0] io_rvfi_regs_30,
  output [63:0] io_rvfi_regs_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [63:0] _RAND_1068;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] PC; // @[cpu.scala 64:19]
  reg [63:0] Regs_0; // @[cpu.scala 65:21]
  reg [63:0] Regs_1; // @[cpu.scala 65:21]
  reg [63:0] Regs_2; // @[cpu.scala 65:21]
  reg [63:0] Regs_3; // @[cpu.scala 65:21]
  reg [63:0] Regs_4; // @[cpu.scala 65:21]
  reg [63:0] Regs_5; // @[cpu.scala 65:21]
  reg [63:0] Regs_6; // @[cpu.scala 65:21]
  reg [63:0] Regs_7; // @[cpu.scala 65:21]
  reg [63:0] Regs_8; // @[cpu.scala 65:21]
  reg [63:0] Regs_9; // @[cpu.scala 65:21]
  reg [63:0] Regs_10; // @[cpu.scala 65:21]
  reg [63:0] Regs_11; // @[cpu.scala 65:21]
  reg [63:0] Regs_12; // @[cpu.scala 65:21]
  reg [63:0] Regs_13; // @[cpu.scala 65:21]
  reg [63:0] Regs_14; // @[cpu.scala 65:21]
  reg [63:0] Regs_15; // @[cpu.scala 65:21]
  reg [63:0] Regs_16; // @[cpu.scala 65:21]
  reg [63:0] Regs_17; // @[cpu.scala 65:21]
  reg [63:0] Regs_18; // @[cpu.scala 65:21]
  reg [63:0] Regs_19; // @[cpu.scala 65:21]
  reg [63:0] Regs_20; // @[cpu.scala 65:21]
  reg [63:0] Regs_21; // @[cpu.scala 65:21]
  reg [63:0] Regs_22; // @[cpu.scala 65:21]
  reg [63:0] Regs_23; // @[cpu.scala 65:21]
  reg [63:0] Regs_24; // @[cpu.scala 65:21]
  reg [63:0] Regs_25; // @[cpu.scala 65:21]
  reg [63:0] Regs_26; // @[cpu.scala 65:21]
  reg [63:0] Regs_27; // @[cpu.scala 65:21]
  reg [63:0] Regs_28; // @[cpu.scala 65:21]
  reg [63:0] Regs_29; // @[cpu.scala 65:21]
  reg [63:0] Regs_30; // @[cpu.scala 65:21]
  reg [63:0] Regs_31; // @[cpu.scala 65:21]
  reg [63:0] IDEXA; // @[cpu.scala 67:58]
  reg [63:0] IDEXB; // @[cpu.scala 67:58]
  reg [63:0] EXMEMB; // @[cpu.scala 67:58]
  reg [63:0] EXMEMALUOut; // @[cpu.scala 67:58]
  reg [63:0] MEMWBValue; // @[cpu.scala 67:58]
  reg [31:0] DMemory_0; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1; // @[cpu.scala 69:24]
  reg [31:0] DMemory_2; // @[cpu.scala 69:24]
  reg [31:0] DMemory_3; // @[cpu.scala 69:24]
  reg [31:0] DMemory_4; // @[cpu.scala 69:24]
  reg [31:0] DMemory_5; // @[cpu.scala 69:24]
  reg [31:0] DMemory_6; // @[cpu.scala 69:24]
  reg [31:0] DMemory_7; // @[cpu.scala 69:24]
  reg [31:0] DMemory_8; // @[cpu.scala 69:24]
  reg [31:0] DMemory_9; // @[cpu.scala 69:24]
  reg [31:0] DMemory_10; // @[cpu.scala 69:24]
  reg [31:0] DMemory_11; // @[cpu.scala 69:24]
  reg [31:0] DMemory_12; // @[cpu.scala 69:24]
  reg [31:0] DMemory_13; // @[cpu.scala 69:24]
  reg [31:0] DMemory_14; // @[cpu.scala 69:24]
  reg [31:0] DMemory_15; // @[cpu.scala 69:24]
  reg [31:0] DMemory_16; // @[cpu.scala 69:24]
  reg [31:0] DMemory_17; // @[cpu.scala 69:24]
  reg [31:0] DMemory_18; // @[cpu.scala 69:24]
  reg [31:0] DMemory_19; // @[cpu.scala 69:24]
  reg [31:0] DMemory_20; // @[cpu.scala 69:24]
  reg [31:0] DMemory_21; // @[cpu.scala 69:24]
  reg [31:0] DMemory_22; // @[cpu.scala 69:24]
  reg [31:0] DMemory_23; // @[cpu.scala 69:24]
  reg [31:0] DMemory_24; // @[cpu.scala 69:24]
  reg [31:0] DMemory_25; // @[cpu.scala 69:24]
  reg [31:0] DMemory_26; // @[cpu.scala 69:24]
  reg [31:0] DMemory_27; // @[cpu.scala 69:24]
  reg [31:0] DMemory_28; // @[cpu.scala 69:24]
  reg [31:0] DMemory_29; // @[cpu.scala 69:24]
  reg [31:0] DMemory_30; // @[cpu.scala 69:24]
  reg [31:0] DMemory_31; // @[cpu.scala 69:24]
  reg [31:0] DMemory_32; // @[cpu.scala 69:24]
  reg [31:0] DMemory_33; // @[cpu.scala 69:24]
  reg [31:0] DMemory_34; // @[cpu.scala 69:24]
  reg [31:0] DMemory_35; // @[cpu.scala 69:24]
  reg [31:0] DMemory_36; // @[cpu.scala 69:24]
  reg [31:0] DMemory_37; // @[cpu.scala 69:24]
  reg [31:0] DMemory_38; // @[cpu.scala 69:24]
  reg [31:0] DMemory_39; // @[cpu.scala 69:24]
  reg [31:0] DMemory_40; // @[cpu.scala 69:24]
  reg [31:0] DMemory_41; // @[cpu.scala 69:24]
  reg [31:0] DMemory_42; // @[cpu.scala 69:24]
  reg [31:0] DMemory_43; // @[cpu.scala 69:24]
  reg [31:0] DMemory_44; // @[cpu.scala 69:24]
  reg [31:0] DMemory_45; // @[cpu.scala 69:24]
  reg [31:0] DMemory_46; // @[cpu.scala 69:24]
  reg [31:0] DMemory_47; // @[cpu.scala 69:24]
  reg [31:0] DMemory_48; // @[cpu.scala 69:24]
  reg [31:0] DMemory_49; // @[cpu.scala 69:24]
  reg [31:0] DMemory_50; // @[cpu.scala 69:24]
  reg [31:0] DMemory_51; // @[cpu.scala 69:24]
  reg [31:0] DMemory_52; // @[cpu.scala 69:24]
  reg [31:0] DMemory_53; // @[cpu.scala 69:24]
  reg [31:0] DMemory_54; // @[cpu.scala 69:24]
  reg [31:0] DMemory_55; // @[cpu.scala 69:24]
  reg [31:0] DMemory_56; // @[cpu.scala 69:24]
  reg [31:0] DMemory_57; // @[cpu.scala 69:24]
  reg [31:0] DMemory_58; // @[cpu.scala 69:24]
  reg [31:0] DMemory_59; // @[cpu.scala 69:24]
  reg [31:0] DMemory_60; // @[cpu.scala 69:24]
  reg [31:0] DMemory_61; // @[cpu.scala 69:24]
  reg [31:0] DMemory_62; // @[cpu.scala 69:24]
  reg [31:0] DMemory_63; // @[cpu.scala 69:24]
  reg [31:0] DMemory_64; // @[cpu.scala 69:24]
  reg [31:0] DMemory_65; // @[cpu.scala 69:24]
  reg [31:0] DMemory_66; // @[cpu.scala 69:24]
  reg [31:0] DMemory_67; // @[cpu.scala 69:24]
  reg [31:0] DMemory_68; // @[cpu.scala 69:24]
  reg [31:0] DMemory_69; // @[cpu.scala 69:24]
  reg [31:0] DMemory_70; // @[cpu.scala 69:24]
  reg [31:0] DMemory_71; // @[cpu.scala 69:24]
  reg [31:0] DMemory_72; // @[cpu.scala 69:24]
  reg [31:0] DMemory_73; // @[cpu.scala 69:24]
  reg [31:0] DMemory_74; // @[cpu.scala 69:24]
  reg [31:0] DMemory_75; // @[cpu.scala 69:24]
  reg [31:0] DMemory_76; // @[cpu.scala 69:24]
  reg [31:0] DMemory_77; // @[cpu.scala 69:24]
  reg [31:0] DMemory_78; // @[cpu.scala 69:24]
  reg [31:0] DMemory_79; // @[cpu.scala 69:24]
  reg [31:0] DMemory_80; // @[cpu.scala 69:24]
  reg [31:0] DMemory_81; // @[cpu.scala 69:24]
  reg [31:0] DMemory_82; // @[cpu.scala 69:24]
  reg [31:0] DMemory_83; // @[cpu.scala 69:24]
  reg [31:0] DMemory_84; // @[cpu.scala 69:24]
  reg [31:0] DMemory_85; // @[cpu.scala 69:24]
  reg [31:0] DMemory_86; // @[cpu.scala 69:24]
  reg [31:0] DMemory_87; // @[cpu.scala 69:24]
  reg [31:0] DMemory_88; // @[cpu.scala 69:24]
  reg [31:0] DMemory_89; // @[cpu.scala 69:24]
  reg [31:0] DMemory_90; // @[cpu.scala 69:24]
  reg [31:0] DMemory_91; // @[cpu.scala 69:24]
  reg [31:0] DMemory_92; // @[cpu.scala 69:24]
  reg [31:0] DMemory_93; // @[cpu.scala 69:24]
  reg [31:0] DMemory_94; // @[cpu.scala 69:24]
  reg [31:0] DMemory_95; // @[cpu.scala 69:24]
  reg [31:0] DMemory_96; // @[cpu.scala 69:24]
  reg [31:0] DMemory_97; // @[cpu.scala 69:24]
  reg [31:0] DMemory_98; // @[cpu.scala 69:24]
  reg [31:0] DMemory_99; // @[cpu.scala 69:24]
  reg [31:0] DMemory_100; // @[cpu.scala 69:24]
  reg [31:0] DMemory_101; // @[cpu.scala 69:24]
  reg [31:0] DMemory_102; // @[cpu.scala 69:24]
  reg [31:0] DMemory_103; // @[cpu.scala 69:24]
  reg [31:0] DMemory_104; // @[cpu.scala 69:24]
  reg [31:0] DMemory_105; // @[cpu.scala 69:24]
  reg [31:0] DMemory_106; // @[cpu.scala 69:24]
  reg [31:0] DMemory_107; // @[cpu.scala 69:24]
  reg [31:0] DMemory_108; // @[cpu.scala 69:24]
  reg [31:0] DMemory_109; // @[cpu.scala 69:24]
  reg [31:0] DMemory_110; // @[cpu.scala 69:24]
  reg [31:0] DMemory_111; // @[cpu.scala 69:24]
  reg [31:0] DMemory_112; // @[cpu.scala 69:24]
  reg [31:0] DMemory_113; // @[cpu.scala 69:24]
  reg [31:0] DMemory_114; // @[cpu.scala 69:24]
  reg [31:0] DMemory_115; // @[cpu.scala 69:24]
  reg [31:0] DMemory_116; // @[cpu.scala 69:24]
  reg [31:0] DMemory_117; // @[cpu.scala 69:24]
  reg [31:0] DMemory_118; // @[cpu.scala 69:24]
  reg [31:0] DMemory_119; // @[cpu.scala 69:24]
  reg [31:0] DMemory_120; // @[cpu.scala 69:24]
  reg [31:0] DMemory_121; // @[cpu.scala 69:24]
  reg [31:0] DMemory_122; // @[cpu.scala 69:24]
  reg [31:0] DMemory_123; // @[cpu.scala 69:24]
  reg [31:0] DMemory_124; // @[cpu.scala 69:24]
  reg [31:0] DMemory_125; // @[cpu.scala 69:24]
  reg [31:0] DMemory_126; // @[cpu.scala 69:24]
  reg [31:0] DMemory_127; // @[cpu.scala 69:24]
  reg [31:0] DMemory_128; // @[cpu.scala 69:24]
  reg [31:0] DMemory_129; // @[cpu.scala 69:24]
  reg [31:0] DMemory_130; // @[cpu.scala 69:24]
  reg [31:0] DMemory_131; // @[cpu.scala 69:24]
  reg [31:0] DMemory_132; // @[cpu.scala 69:24]
  reg [31:0] DMemory_133; // @[cpu.scala 69:24]
  reg [31:0] DMemory_134; // @[cpu.scala 69:24]
  reg [31:0] DMemory_135; // @[cpu.scala 69:24]
  reg [31:0] DMemory_136; // @[cpu.scala 69:24]
  reg [31:0] DMemory_137; // @[cpu.scala 69:24]
  reg [31:0] DMemory_138; // @[cpu.scala 69:24]
  reg [31:0] DMemory_139; // @[cpu.scala 69:24]
  reg [31:0] DMemory_140; // @[cpu.scala 69:24]
  reg [31:0] DMemory_141; // @[cpu.scala 69:24]
  reg [31:0] DMemory_142; // @[cpu.scala 69:24]
  reg [31:0] DMemory_143; // @[cpu.scala 69:24]
  reg [31:0] DMemory_144; // @[cpu.scala 69:24]
  reg [31:0] DMemory_145; // @[cpu.scala 69:24]
  reg [31:0] DMemory_146; // @[cpu.scala 69:24]
  reg [31:0] DMemory_147; // @[cpu.scala 69:24]
  reg [31:0] DMemory_148; // @[cpu.scala 69:24]
  reg [31:0] DMemory_149; // @[cpu.scala 69:24]
  reg [31:0] DMemory_150; // @[cpu.scala 69:24]
  reg [31:0] DMemory_151; // @[cpu.scala 69:24]
  reg [31:0] DMemory_152; // @[cpu.scala 69:24]
  reg [31:0] DMemory_153; // @[cpu.scala 69:24]
  reg [31:0] DMemory_154; // @[cpu.scala 69:24]
  reg [31:0] DMemory_155; // @[cpu.scala 69:24]
  reg [31:0] DMemory_156; // @[cpu.scala 69:24]
  reg [31:0] DMemory_157; // @[cpu.scala 69:24]
  reg [31:0] DMemory_158; // @[cpu.scala 69:24]
  reg [31:0] DMemory_159; // @[cpu.scala 69:24]
  reg [31:0] DMemory_160; // @[cpu.scala 69:24]
  reg [31:0] DMemory_161; // @[cpu.scala 69:24]
  reg [31:0] DMemory_162; // @[cpu.scala 69:24]
  reg [31:0] DMemory_163; // @[cpu.scala 69:24]
  reg [31:0] DMemory_164; // @[cpu.scala 69:24]
  reg [31:0] DMemory_165; // @[cpu.scala 69:24]
  reg [31:0] DMemory_166; // @[cpu.scala 69:24]
  reg [31:0] DMemory_167; // @[cpu.scala 69:24]
  reg [31:0] DMemory_168; // @[cpu.scala 69:24]
  reg [31:0] DMemory_169; // @[cpu.scala 69:24]
  reg [31:0] DMemory_170; // @[cpu.scala 69:24]
  reg [31:0] DMemory_171; // @[cpu.scala 69:24]
  reg [31:0] DMemory_172; // @[cpu.scala 69:24]
  reg [31:0] DMemory_173; // @[cpu.scala 69:24]
  reg [31:0] DMemory_174; // @[cpu.scala 69:24]
  reg [31:0] DMemory_175; // @[cpu.scala 69:24]
  reg [31:0] DMemory_176; // @[cpu.scala 69:24]
  reg [31:0] DMemory_177; // @[cpu.scala 69:24]
  reg [31:0] DMemory_178; // @[cpu.scala 69:24]
  reg [31:0] DMemory_179; // @[cpu.scala 69:24]
  reg [31:0] DMemory_180; // @[cpu.scala 69:24]
  reg [31:0] DMemory_181; // @[cpu.scala 69:24]
  reg [31:0] DMemory_182; // @[cpu.scala 69:24]
  reg [31:0] DMemory_183; // @[cpu.scala 69:24]
  reg [31:0] DMemory_184; // @[cpu.scala 69:24]
  reg [31:0] DMemory_185; // @[cpu.scala 69:24]
  reg [31:0] DMemory_186; // @[cpu.scala 69:24]
  reg [31:0] DMemory_187; // @[cpu.scala 69:24]
  reg [31:0] DMemory_188; // @[cpu.scala 69:24]
  reg [31:0] DMemory_189; // @[cpu.scala 69:24]
  reg [31:0] DMemory_190; // @[cpu.scala 69:24]
  reg [31:0] DMemory_191; // @[cpu.scala 69:24]
  reg [31:0] DMemory_192; // @[cpu.scala 69:24]
  reg [31:0] DMemory_193; // @[cpu.scala 69:24]
  reg [31:0] DMemory_194; // @[cpu.scala 69:24]
  reg [31:0] DMemory_195; // @[cpu.scala 69:24]
  reg [31:0] DMemory_196; // @[cpu.scala 69:24]
  reg [31:0] DMemory_197; // @[cpu.scala 69:24]
  reg [31:0] DMemory_198; // @[cpu.scala 69:24]
  reg [31:0] DMemory_199; // @[cpu.scala 69:24]
  reg [31:0] DMemory_200; // @[cpu.scala 69:24]
  reg [31:0] DMemory_201; // @[cpu.scala 69:24]
  reg [31:0] DMemory_202; // @[cpu.scala 69:24]
  reg [31:0] DMemory_203; // @[cpu.scala 69:24]
  reg [31:0] DMemory_204; // @[cpu.scala 69:24]
  reg [31:0] DMemory_205; // @[cpu.scala 69:24]
  reg [31:0] DMemory_206; // @[cpu.scala 69:24]
  reg [31:0] DMemory_207; // @[cpu.scala 69:24]
  reg [31:0] DMemory_208; // @[cpu.scala 69:24]
  reg [31:0] DMemory_209; // @[cpu.scala 69:24]
  reg [31:0] DMemory_210; // @[cpu.scala 69:24]
  reg [31:0] DMemory_211; // @[cpu.scala 69:24]
  reg [31:0] DMemory_212; // @[cpu.scala 69:24]
  reg [31:0] DMemory_213; // @[cpu.scala 69:24]
  reg [31:0] DMemory_214; // @[cpu.scala 69:24]
  reg [31:0] DMemory_215; // @[cpu.scala 69:24]
  reg [31:0] DMemory_216; // @[cpu.scala 69:24]
  reg [31:0] DMemory_217; // @[cpu.scala 69:24]
  reg [31:0] DMemory_218; // @[cpu.scala 69:24]
  reg [31:0] DMemory_219; // @[cpu.scala 69:24]
  reg [31:0] DMemory_220; // @[cpu.scala 69:24]
  reg [31:0] DMemory_221; // @[cpu.scala 69:24]
  reg [31:0] DMemory_222; // @[cpu.scala 69:24]
  reg [31:0] DMemory_223; // @[cpu.scala 69:24]
  reg [31:0] DMemory_224; // @[cpu.scala 69:24]
  reg [31:0] DMemory_225; // @[cpu.scala 69:24]
  reg [31:0] DMemory_226; // @[cpu.scala 69:24]
  reg [31:0] DMemory_227; // @[cpu.scala 69:24]
  reg [31:0] DMemory_228; // @[cpu.scala 69:24]
  reg [31:0] DMemory_229; // @[cpu.scala 69:24]
  reg [31:0] DMemory_230; // @[cpu.scala 69:24]
  reg [31:0] DMemory_231; // @[cpu.scala 69:24]
  reg [31:0] DMemory_232; // @[cpu.scala 69:24]
  reg [31:0] DMemory_233; // @[cpu.scala 69:24]
  reg [31:0] DMemory_234; // @[cpu.scala 69:24]
  reg [31:0] DMemory_235; // @[cpu.scala 69:24]
  reg [31:0] DMemory_236; // @[cpu.scala 69:24]
  reg [31:0] DMemory_237; // @[cpu.scala 69:24]
  reg [31:0] DMemory_238; // @[cpu.scala 69:24]
  reg [31:0] DMemory_239; // @[cpu.scala 69:24]
  reg [31:0] DMemory_240; // @[cpu.scala 69:24]
  reg [31:0] DMemory_241; // @[cpu.scala 69:24]
  reg [31:0] DMemory_242; // @[cpu.scala 69:24]
  reg [31:0] DMemory_243; // @[cpu.scala 69:24]
  reg [31:0] DMemory_244; // @[cpu.scala 69:24]
  reg [31:0] DMemory_245; // @[cpu.scala 69:24]
  reg [31:0] DMemory_246; // @[cpu.scala 69:24]
  reg [31:0] DMemory_247; // @[cpu.scala 69:24]
  reg [31:0] DMemory_248; // @[cpu.scala 69:24]
  reg [31:0] DMemory_249; // @[cpu.scala 69:24]
  reg [31:0] DMemory_250; // @[cpu.scala 69:24]
  reg [31:0] DMemory_251; // @[cpu.scala 69:24]
  reg [31:0] DMemory_252; // @[cpu.scala 69:24]
  reg [31:0] DMemory_253; // @[cpu.scala 69:24]
  reg [31:0] DMemory_254; // @[cpu.scala 69:24]
  reg [31:0] DMemory_255; // @[cpu.scala 69:24]
  reg [31:0] DMemory_256; // @[cpu.scala 69:24]
  reg [31:0] DMemory_257; // @[cpu.scala 69:24]
  reg [31:0] DMemory_258; // @[cpu.scala 69:24]
  reg [31:0] DMemory_259; // @[cpu.scala 69:24]
  reg [31:0] DMemory_260; // @[cpu.scala 69:24]
  reg [31:0] DMemory_261; // @[cpu.scala 69:24]
  reg [31:0] DMemory_262; // @[cpu.scala 69:24]
  reg [31:0] DMemory_263; // @[cpu.scala 69:24]
  reg [31:0] DMemory_264; // @[cpu.scala 69:24]
  reg [31:0] DMemory_265; // @[cpu.scala 69:24]
  reg [31:0] DMemory_266; // @[cpu.scala 69:24]
  reg [31:0] DMemory_267; // @[cpu.scala 69:24]
  reg [31:0] DMemory_268; // @[cpu.scala 69:24]
  reg [31:0] DMemory_269; // @[cpu.scala 69:24]
  reg [31:0] DMemory_270; // @[cpu.scala 69:24]
  reg [31:0] DMemory_271; // @[cpu.scala 69:24]
  reg [31:0] DMemory_272; // @[cpu.scala 69:24]
  reg [31:0] DMemory_273; // @[cpu.scala 69:24]
  reg [31:0] DMemory_274; // @[cpu.scala 69:24]
  reg [31:0] DMemory_275; // @[cpu.scala 69:24]
  reg [31:0] DMemory_276; // @[cpu.scala 69:24]
  reg [31:0] DMemory_277; // @[cpu.scala 69:24]
  reg [31:0] DMemory_278; // @[cpu.scala 69:24]
  reg [31:0] DMemory_279; // @[cpu.scala 69:24]
  reg [31:0] DMemory_280; // @[cpu.scala 69:24]
  reg [31:0] DMemory_281; // @[cpu.scala 69:24]
  reg [31:0] DMemory_282; // @[cpu.scala 69:24]
  reg [31:0] DMemory_283; // @[cpu.scala 69:24]
  reg [31:0] DMemory_284; // @[cpu.scala 69:24]
  reg [31:0] DMemory_285; // @[cpu.scala 69:24]
  reg [31:0] DMemory_286; // @[cpu.scala 69:24]
  reg [31:0] DMemory_287; // @[cpu.scala 69:24]
  reg [31:0] DMemory_288; // @[cpu.scala 69:24]
  reg [31:0] DMemory_289; // @[cpu.scala 69:24]
  reg [31:0] DMemory_290; // @[cpu.scala 69:24]
  reg [31:0] DMemory_291; // @[cpu.scala 69:24]
  reg [31:0] DMemory_292; // @[cpu.scala 69:24]
  reg [31:0] DMemory_293; // @[cpu.scala 69:24]
  reg [31:0] DMemory_294; // @[cpu.scala 69:24]
  reg [31:0] DMemory_295; // @[cpu.scala 69:24]
  reg [31:0] DMemory_296; // @[cpu.scala 69:24]
  reg [31:0] DMemory_297; // @[cpu.scala 69:24]
  reg [31:0] DMemory_298; // @[cpu.scala 69:24]
  reg [31:0] DMemory_299; // @[cpu.scala 69:24]
  reg [31:0] DMemory_300; // @[cpu.scala 69:24]
  reg [31:0] DMemory_301; // @[cpu.scala 69:24]
  reg [31:0] DMemory_302; // @[cpu.scala 69:24]
  reg [31:0] DMemory_303; // @[cpu.scala 69:24]
  reg [31:0] DMemory_304; // @[cpu.scala 69:24]
  reg [31:0] DMemory_305; // @[cpu.scala 69:24]
  reg [31:0] DMemory_306; // @[cpu.scala 69:24]
  reg [31:0] DMemory_307; // @[cpu.scala 69:24]
  reg [31:0] DMemory_308; // @[cpu.scala 69:24]
  reg [31:0] DMemory_309; // @[cpu.scala 69:24]
  reg [31:0] DMemory_310; // @[cpu.scala 69:24]
  reg [31:0] DMemory_311; // @[cpu.scala 69:24]
  reg [31:0] DMemory_312; // @[cpu.scala 69:24]
  reg [31:0] DMemory_313; // @[cpu.scala 69:24]
  reg [31:0] DMemory_314; // @[cpu.scala 69:24]
  reg [31:0] DMemory_315; // @[cpu.scala 69:24]
  reg [31:0] DMemory_316; // @[cpu.scala 69:24]
  reg [31:0] DMemory_317; // @[cpu.scala 69:24]
  reg [31:0] DMemory_318; // @[cpu.scala 69:24]
  reg [31:0] DMemory_319; // @[cpu.scala 69:24]
  reg [31:0] DMemory_320; // @[cpu.scala 69:24]
  reg [31:0] DMemory_321; // @[cpu.scala 69:24]
  reg [31:0] DMemory_322; // @[cpu.scala 69:24]
  reg [31:0] DMemory_323; // @[cpu.scala 69:24]
  reg [31:0] DMemory_324; // @[cpu.scala 69:24]
  reg [31:0] DMemory_325; // @[cpu.scala 69:24]
  reg [31:0] DMemory_326; // @[cpu.scala 69:24]
  reg [31:0] DMemory_327; // @[cpu.scala 69:24]
  reg [31:0] DMemory_328; // @[cpu.scala 69:24]
  reg [31:0] DMemory_329; // @[cpu.scala 69:24]
  reg [31:0] DMemory_330; // @[cpu.scala 69:24]
  reg [31:0] DMemory_331; // @[cpu.scala 69:24]
  reg [31:0] DMemory_332; // @[cpu.scala 69:24]
  reg [31:0] DMemory_333; // @[cpu.scala 69:24]
  reg [31:0] DMemory_334; // @[cpu.scala 69:24]
  reg [31:0] DMemory_335; // @[cpu.scala 69:24]
  reg [31:0] DMemory_336; // @[cpu.scala 69:24]
  reg [31:0] DMemory_337; // @[cpu.scala 69:24]
  reg [31:0] DMemory_338; // @[cpu.scala 69:24]
  reg [31:0] DMemory_339; // @[cpu.scala 69:24]
  reg [31:0] DMemory_340; // @[cpu.scala 69:24]
  reg [31:0] DMemory_341; // @[cpu.scala 69:24]
  reg [31:0] DMemory_342; // @[cpu.scala 69:24]
  reg [31:0] DMemory_343; // @[cpu.scala 69:24]
  reg [31:0] DMemory_344; // @[cpu.scala 69:24]
  reg [31:0] DMemory_345; // @[cpu.scala 69:24]
  reg [31:0] DMemory_346; // @[cpu.scala 69:24]
  reg [31:0] DMemory_347; // @[cpu.scala 69:24]
  reg [31:0] DMemory_348; // @[cpu.scala 69:24]
  reg [31:0] DMemory_349; // @[cpu.scala 69:24]
  reg [31:0] DMemory_350; // @[cpu.scala 69:24]
  reg [31:0] DMemory_351; // @[cpu.scala 69:24]
  reg [31:0] DMemory_352; // @[cpu.scala 69:24]
  reg [31:0] DMemory_353; // @[cpu.scala 69:24]
  reg [31:0] DMemory_354; // @[cpu.scala 69:24]
  reg [31:0] DMemory_355; // @[cpu.scala 69:24]
  reg [31:0] DMemory_356; // @[cpu.scala 69:24]
  reg [31:0] DMemory_357; // @[cpu.scala 69:24]
  reg [31:0] DMemory_358; // @[cpu.scala 69:24]
  reg [31:0] DMemory_359; // @[cpu.scala 69:24]
  reg [31:0] DMemory_360; // @[cpu.scala 69:24]
  reg [31:0] DMemory_361; // @[cpu.scala 69:24]
  reg [31:0] DMemory_362; // @[cpu.scala 69:24]
  reg [31:0] DMemory_363; // @[cpu.scala 69:24]
  reg [31:0] DMemory_364; // @[cpu.scala 69:24]
  reg [31:0] DMemory_365; // @[cpu.scala 69:24]
  reg [31:0] DMemory_366; // @[cpu.scala 69:24]
  reg [31:0] DMemory_367; // @[cpu.scala 69:24]
  reg [31:0] DMemory_368; // @[cpu.scala 69:24]
  reg [31:0] DMemory_369; // @[cpu.scala 69:24]
  reg [31:0] DMemory_370; // @[cpu.scala 69:24]
  reg [31:0] DMemory_371; // @[cpu.scala 69:24]
  reg [31:0] DMemory_372; // @[cpu.scala 69:24]
  reg [31:0] DMemory_373; // @[cpu.scala 69:24]
  reg [31:0] DMemory_374; // @[cpu.scala 69:24]
  reg [31:0] DMemory_375; // @[cpu.scala 69:24]
  reg [31:0] DMemory_376; // @[cpu.scala 69:24]
  reg [31:0] DMemory_377; // @[cpu.scala 69:24]
  reg [31:0] DMemory_378; // @[cpu.scala 69:24]
  reg [31:0] DMemory_379; // @[cpu.scala 69:24]
  reg [31:0] DMemory_380; // @[cpu.scala 69:24]
  reg [31:0] DMemory_381; // @[cpu.scala 69:24]
  reg [31:0] DMemory_382; // @[cpu.scala 69:24]
  reg [31:0] DMemory_383; // @[cpu.scala 69:24]
  reg [31:0] DMemory_384; // @[cpu.scala 69:24]
  reg [31:0] DMemory_385; // @[cpu.scala 69:24]
  reg [31:0] DMemory_386; // @[cpu.scala 69:24]
  reg [31:0] DMemory_387; // @[cpu.scala 69:24]
  reg [31:0] DMemory_388; // @[cpu.scala 69:24]
  reg [31:0] DMemory_389; // @[cpu.scala 69:24]
  reg [31:0] DMemory_390; // @[cpu.scala 69:24]
  reg [31:0] DMemory_391; // @[cpu.scala 69:24]
  reg [31:0] DMemory_392; // @[cpu.scala 69:24]
  reg [31:0] DMemory_393; // @[cpu.scala 69:24]
  reg [31:0] DMemory_394; // @[cpu.scala 69:24]
  reg [31:0] DMemory_395; // @[cpu.scala 69:24]
  reg [31:0] DMemory_396; // @[cpu.scala 69:24]
  reg [31:0] DMemory_397; // @[cpu.scala 69:24]
  reg [31:0] DMemory_398; // @[cpu.scala 69:24]
  reg [31:0] DMemory_399; // @[cpu.scala 69:24]
  reg [31:0] DMemory_400; // @[cpu.scala 69:24]
  reg [31:0] DMemory_401; // @[cpu.scala 69:24]
  reg [31:0] DMemory_402; // @[cpu.scala 69:24]
  reg [31:0] DMemory_403; // @[cpu.scala 69:24]
  reg [31:0] DMemory_404; // @[cpu.scala 69:24]
  reg [31:0] DMemory_405; // @[cpu.scala 69:24]
  reg [31:0] DMemory_406; // @[cpu.scala 69:24]
  reg [31:0] DMemory_407; // @[cpu.scala 69:24]
  reg [31:0] DMemory_408; // @[cpu.scala 69:24]
  reg [31:0] DMemory_409; // @[cpu.scala 69:24]
  reg [31:0] DMemory_410; // @[cpu.scala 69:24]
  reg [31:0] DMemory_411; // @[cpu.scala 69:24]
  reg [31:0] DMemory_412; // @[cpu.scala 69:24]
  reg [31:0] DMemory_413; // @[cpu.scala 69:24]
  reg [31:0] DMemory_414; // @[cpu.scala 69:24]
  reg [31:0] DMemory_415; // @[cpu.scala 69:24]
  reg [31:0] DMemory_416; // @[cpu.scala 69:24]
  reg [31:0] DMemory_417; // @[cpu.scala 69:24]
  reg [31:0] DMemory_418; // @[cpu.scala 69:24]
  reg [31:0] DMemory_419; // @[cpu.scala 69:24]
  reg [31:0] DMemory_420; // @[cpu.scala 69:24]
  reg [31:0] DMemory_421; // @[cpu.scala 69:24]
  reg [31:0] DMemory_422; // @[cpu.scala 69:24]
  reg [31:0] DMemory_423; // @[cpu.scala 69:24]
  reg [31:0] DMemory_424; // @[cpu.scala 69:24]
  reg [31:0] DMemory_425; // @[cpu.scala 69:24]
  reg [31:0] DMemory_426; // @[cpu.scala 69:24]
  reg [31:0] DMemory_427; // @[cpu.scala 69:24]
  reg [31:0] DMemory_428; // @[cpu.scala 69:24]
  reg [31:0] DMemory_429; // @[cpu.scala 69:24]
  reg [31:0] DMemory_430; // @[cpu.scala 69:24]
  reg [31:0] DMemory_431; // @[cpu.scala 69:24]
  reg [31:0] DMemory_432; // @[cpu.scala 69:24]
  reg [31:0] DMemory_433; // @[cpu.scala 69:24]
  reg [31:0] DMemory_434; // @[cpu.scala 69:24]
  reg [31:0] DMemory_435; // @[cpu.scala 69:24]
  reg [31:0] DMemory_436; // @[cpu.scala 69:24]
  reg [31:0] DMemory_437; // @[cpu.scala 69:24]
  reg [31:0] DMemory_438; // @[cpu.scala 69:24]
  reg [31:0] DMemory_439; // @[cpu.scala 69:24]
  reg [31:0] DMemory_440; // @[cpu.scala 69:24]
  reg [31:0] DMemory_441; // @[cpu.scala 69:24]
  reg [31:0] DMemory_442; // @[cpu.scala 69:24]
  reg [31:0] DMemory_443; // @[cpu.scala 69:24]
  reg [31:0] DMemory_444; // @[cpu.scala 69:24]
  reg [31:0] DMemory_445; // @[cpu.scala 69:24]
  reg [31:0] DMemory_446; // @[cpu.scala 69:24]
  reg [31:0] DMemory_447; // @[cpu.scala 69:24]
  reg [31:0] DMemory_448; // @[cpu.scala 69:24]
  reg [31:0] DMemory_449; // @[cpu.scala 69:24]
  reg [31:0] DMemory_450; // @[cpu.scala 69:24]
  reg [31:0] DMemory_451; // @[cpu.scala 69:24]
  reg [31:0] DMemory_452; // @[cpu.scala 69:24]
  reg [31:0] DMemory_453; // @[cpu.scala 69:24]
  reg [31:0] DMemory_454; // @[cpu.scala 69:24]
  reg [31:0] DMemory_455; // @[cpu.scala 69:24]
  reg [31:0] DMemory_456; // @[cpu.scala 69:24]
  reg [31:0] DMemory_457; // @[cpu.scala 69:24]
  reg [31:0] DMemory_458; // @[cpu.scala 69:24]
  reg [31:0] DMemory_459; // @[cpu.scala 69:24]
  reg [31:0] DMemory_460; // @[cpu.scala 69:24]
  reg [31:0] DMemory_461; // @[cpu.scala 69:24]
  reg [31:0] DMemory_462; // @[cpu.scala 69:24]
  reg [31:0] DMemory_463; // @[cpu.scala 69:24]
  reg [31:0] DMemory_464; // @[cpu.scala 69:24]
  reg [31:0] DMemory_465; // @[cpu.scala 69:24]
  reg [31:0] DMemory_466; // @[cpu.scala 69:24]
  reg [31:0] DMemory_467; // @[cpu.scala 69:24]
  reg [31:0] DMemory_468; // @[cpu.scala 69:24]
  reg [31:0] DMemory_469; // @[cpu.scala 69:24]
  reg [31:0] DMemory_470; // @[cpu.scala 69:24]
  reg [31:0] DMemory_471; // @[cpu.scala 69:24]
  reg [31:0] DMemory_472; // @[cpu.scala 69:24]
  reg [31:0] DMemory_473; // @[cpu.scala 69:24]
  reg [31:0] DMemory_474; // @[cpu.scala 69:24]
  reg [31:0] DMemory_475; // @[cpu.scala 69:24]
  reg [31:0] DMemory_476; // @[cpu.scala 69:24]
  reg [31:0] DMemory_477; // @[cpu.scala 69:24]
  reg [31:0] DMemory_478; // @[cpu.scala 69:24]
  reg [31:0] DMemory_479; // @[cpu.scala 69:24]
  reg [31:0] DMemory_480; // @[cpu.scala 69:24]
  reg [31:0] DMemory_481; // @[cpu.scala 69:24]
  reg [31:0] DMemory_482; // @[cpu.scala 69:24]
  reg [31:0] DMemory_483; // @[cpu.scala 69:24]
  reg [31:0] DMemory_484; // @[cpu.scala 69:24]
  reg [31:0] DMemory_485; // @[cpu.scala 69:24]
  reg [31:0] DMemory_486; // @[cpu.scala 69:24]
  reg [31:0] DMemory_487; // @[cpu.scala 69:24]
  reg [31:0] DMemory_488; // @[cpu.scala 69:24]
  reg [31:0] DMemory_489; // @[cpu.scala 69:24]
  reg [31:0] DMemory_490; // @[cpu.scala 69:24]
  reg [31:0] DMemory_491; // @[cpu.scala 69:24]
  reg [31:0] DMemory_492; // @[cpu.scala 69:24]
  reg [31:0] DMemory_493; // @[cpu.scala 69:24]
  reg [31:0] DMemory_494; // @[cpu.scala 69:24]
  reg [31:0] DMemory_495; // @[cpu.scala 69:24]
  reg [31:0] DMemory_496; // @[cpu.scala 69:24]
  reg [31:0] DMemory_497; // @[cpu.scala 69:24]
  reg [31:0] DMemory_498; // @[cpu.scala 69:24]
  reg [31:0] DMemory_499; // @[cpu.scala 69:24]
  reg [31:0] DMemory_500; // @[cpu.scala 69:24]
  reg [31:0] DMemory_501; // @[cpu.scala 69:24]
  reg [31:0] DMemory_502; // @[cpu.scala 69:24]
  reg [31:0] DMemory_503; // @[cpu.scala 69:24]
  reg [31:0] DMemory_504; // @[cpu.scala 69:24]
  reg [31:0] DMemory_505; // @[cpu.scala 69:24]
  reg [31:0] DMemory_506; // @[cpu.scala 69:24]
  reg [31:0] DMemory_507; // @[cpu.scala 69:24]
  reg [31:0] DMemory_508; // @[cpu.scala 69:24]
  reg [31:0] DMemory_509; // @[cpu.scala 69:24]
  reg [31:0] DMemory_510; // @[cpu.scala 69:24]
  reg [31:0] DMemory_511; // @[cpu.scala 69:24]
  reg [31:0] DMemory_512; // @[cpu.scala 69:24]
  reg [31:0] DMemory_513; // @[cpu.scala 69:24]
  reg [31:0] DMemory_514; // @[cpu.scala 69:24]
  reg [31:0] DMemory_515; // @[cpu.scala 69:24]
  reg [31:0] DMemory_516; // @[cpu.scala 69:24]
  reg [31:0] DMemory_517; // @[cpu.scala 69:24]
  reg [31:0] DMemory_518; // @[cpu.scala 69:24]
  reg [31:0] DMemory_519; // @[cpu.scala 69:24]
  reg [31:0] DMemory_520; // @[cpu.scala 69:24]
  reg [31:0] DMemory_521; // @[cpu.scala 69:24]
  reg [31:0] DMemory_522; // @[cpu.scala 69:24]
  reg [31:0] DMemory_523; // @[cpu.scala 69:24]
  reg [31:0] DMemory_524; // @[cpu.scala 69:24]
  reg [31:0] DMemory_525; // @[cpu.scala 69:24]
  reg [31:0] DMemory_526; // @[cpu.scala 69:24]
  reg [31:0] DMemory_527; // @[cpu.scala 69:24]
  reg [31:0] DMemory_528; // @[cpu.scala 69:24]
  reg [31:0] DMemory_529; // @[cpu.scala 69:24]
  reg [31:0] DMemory_530; // @[cpu.scala 69:24]
  reg [31:0] DMemory_531; // @[cpu.scala 69:24]
  reg [31:0] DMemory_532; // @[cpu.scala 69:24]
  reg [31:0] DMemory_533; // @[cpu.scala 69:24]
  reg [31:0] DMemory_534; // @[cpu.scala 69:24]
  reg [31:0] DMemory_535; // @[cpu.scala 69:24]
  reg [31:0] DMemory_536; // @[cpu.scala 69:24]
  reg [31:0] DMemory_537; // @[cpu.scala 69:24]
  reg [31:0] DMemory_538; // @[cpu.scala 69:24]
  reg [31:0] DMemory_539; // @[cpu.scala 69:24]
  reg [31:0] DMemory_540; // @[cpu.scala 69:24]
  reg [31:0] DMemory_541; // @[cpu.scala 69:24]
  reg [31:0] DMemory_542; // @[cpu.scala 69:24]
  reg [31:0] DMemory_543; // @[cpu.scala 69:24]
  reg [31:0] DMemory_544; // @[cpu.scala 69:24]
  reg [31:0] DMemory_545; // @[cpu.scala 69:24]
  reg [31:0] DMemory_546; // @[cpu.scala 69:24]
  reg [31:0] DMemory_547; // @[cpu.scala 69:24]
  reg [31:0] DMemory_548; // @[cpu.scala 69:24]
  reg [31:0] DMemory_549; // @[cpu.scala 69:24]
  reg [31:0] DMemory_550; // @[cpu.scala 69:24]
  reg [31:0] DMemory_551; // @[cpu.scala 69:24]
  reg [31:0] DMemory_552; // @[cpu.scala 69:24]
  reg [31:0] DMemory_553; // @[cpu.scala 69:24]
  reg [31:0] DMemory_554; // @[cpu.scala 69:24]
  reg [31:0] DMemory_555; // @[cpu.scala 69:24]
  reg [31:0] DMemory_556; // @[cpu.scala 69:24]
  reg [31:0] DMemory_557; // @[cpu.scala 69:24]
  reg [31:0] DMemory_558; // @[cpu.scala 69:24]
  reg [31:0] DMemory_559; // @[cpu.scala 69:24]
  reg [31:0] DMemory_560; // @[cpu.scala 69:24]
  reg [31:0] DMemory_561; // @[cpu.scala 69:24]
  reg [31:0] DMemory_562; // @[cpu.scala 69:24]
  reg [31:0] DMemory_563; // @[cpu.scala 69:24]
  reg [31:0] DMemory_564; // @[cpu.scala 69:24]
  reg [31:0] DMemory_565; // @[cpu.scala 69:24]
  reg [31:0] DMemory_566; // @[cpu.scala 69:24]
  reg [31:0] DMemory_567; // @[cpu.scala 69:24]
  reg [31:0] DMemory_568; // @[cpu.scala 69:24]
  reg [31:0] DMemory_569; // @[cpu.scala 69:24]
  reg [31:0] DMemory_570; // @[cpu.scala 69:24]
  reg [31:0] DMemory_571; // @[cpu.scala 69:24]
  reg [31:0] DMemory_572; // @[cpu.scala 69:24]
  reg [31:0] DMemory_573; // @[cpu.scala 69:24]
  reg [31:0] DMemory_574; // @[cpu.scala 69:24]
  reg [31:0] DMemory_575; // @[cpu.scala 69:24]
  reg [31:0] DMemory_576; // @[cpu.scala 69:24]
  reg [31:0] DMemory_577; // @[cpu.scala 69:24]
  reg [31:0] DMemory_578; // @[cpu.scala 69:24]
  reg [31:0] DMemory_579; // @[cpu.scala 69:24]
  reg [31:0] DMemory_580; // @[cpu.scala 69:24]
  reg [31:0] DMemory_581; // @[cpu.scala 69:24]
  reg [31:0] DMemory_582; // @[cpu.scala 69:24]
  reg [31:0] DMemory_583; // @[cpu.scala 69:24]
  reg [31:0] DMemory_584; // @[cpu.scala 69:24]
  reg [31:0] DMemory_585; // @[cpu.scala 69:24]
  reg [31:0] DMemory_586; // @[cpu.scala 69:24]
  reg [31:0] DMemory_587; // @[cpu.scala 69:24]
  reg [31:0] DMemory_588; // @[cpu.scala 69:24]
  reg [31:0] DMemory_589; // @[cpu.scala 69:24]
  reg [31:0] DMemory_590; // @[cpu.scala 69:24]
  reg [31:0] DMemory_591; // @[cpu.scala 69:24]
  reg [31:0] DMemory_592; // @[cpu.scala 69:24]
  reg [31:0] DMemory_593; // @[cpu.scala 69:24]
  reg [31:0] DMemory_594; // @[cpu.scala 69:24]
  reg [31:0] DMemory_595; // @[cpu.scala 69:24]
  reg [31:0] DMemory_596; // @[cpu.scala 69:24]
  reg [31:0] DMemory_597; // @[cpu.scala 69:24]
  reg [31:0] DMemory_598; // @[cpu.scala 69:24]
  reg [31:0] DMemory_599; // @[cpu.scala 69:24]
  reg [31:0] DMemory_600; // @[cpu.scala 69:24]
  reg [31:0] DMemory_601; // @[cpu.scala 69:24]
  reg [31:0] DMemory_602; // @[cpu.scala 69:24]
  reg [31:0] DMemory_603; // @[cpu.scala 69:24]
  reg [31:0] DMemory_604; // @[cpu.scala 69:24]
  reg [31:0] DMemory_605; // @[cpu.scala 69:24]
  reg [31:0] DMemory_606; // @[cpu.scala 69:24]
  reg [31:0] DMemory_607; // @[cpu.scala 69:24]
  reg [31:0] DMemory_608; // @[cpu.scala 69:24]
  reg [31:0] DMemory_609; // @[cpu.scala 69:24]
  reg [31:0] DMemory_610; // @[cpu.scala 69:24]
  reg [31:0] DMemory_611; // @[cpu.scala 69:24]
  reg [31:0] DMemory_612; // @[cpu.scala 69:24]
  reg [31:0] DMemory_613; // @[cpu.scala 69:24]
  reg [31:0] DMemory_614; // @[cpu.scala 69:24]
  reg [31:0] DMemory_615; // @[cpu.scala 69:24]
  reg [31:0] DMemory_616; // @[cpu.scala 69:24]
  reg [31:0] DMemory_617; // @[cpu.scala 69:24]
  reg [31:0] DMemory_618; // @[cpu.scala 69:24]
  reg [31:0] DMemory_619; // @[cpu.scala 69:24]
  reg [31:0] DMemory_620; // @[cpu.scala 69:24]
  reg [31:0] DMemory_621; // @[cpu.scala 69:24]
  reg [31:0] DMemory_622; // @[cpu.scala 69:24]
  reg [31:0] DMemory_623; // @[cpu.scala 69:24]
  reg [31:0] DMemory_624; // @[cpu.scala 69:24]
  reg [31:0] DMemory_625; // @[cpu.scala 69:24]
  reg [31:0] DMemory_626; // @[cpu.scala 69:24]
  reg [31:0] DMemory_627; // @[cpu.scala 69:24]
  reg [31:0] DMemory_628; // @[cpu.scala 69:24]
  reg [31:0] DMemory_629; // @[cpu.scala 69:24]
  reg [31:0] DMemory_630; // @[cpu.scala 69:24]
  reg [31:0] DMemory_631; // @[cpu.scala 69:24]
  reg [31:0] DMemory_632; // @[cpu.scala 69:24]
  reg [31:0] DMemory_633; // @[cpu.scala 69:24]
  reg [31:0] DMemory_634; // @[cpu.scala 69:24]
  reg [31:0] DMemory_635; // @[cpu.scala 69:24]
  reg [31:0] DMemory_636; // @[cpu.scala 69:24]
  reg [31:0] DMemory_637; // @[cpu.scala 69:24]
  reg [31:0] DMemory_638; // @[cpu.scala 69:24]
  reg [31:0] DMemory_639; // @[cpu.scala 69:24]
  reg [31:0] DMemory_640; // @[cpu.scala 69:24]
  reg [31:0] DMemory_641; // @[cpu.scala 69:24]
  reg [31:0] DMemory_642; // @[cpu.scala 69:24]
  reg [31:0] DMemory_643; // @[cpu.scala 69:24]
  reg [31:0] DMemory_644; // @[cpu.scala 69:24]
  reg [31:0] DMemory_645; // @[cpu.scala 69:24]
  reg [31:0] DMemory_646; // @[cpu.scala 69:24]
  reg [31:0] DMemory_647; // @[cpu.scala 69:24]
  reg [31:0] DMemory_648; // @[cpu.scala 69:24]
  reg [31:0] DMemory_649; // @[cpu.scala 69:24]
  reg [31:0] DMemory_650; // @[cpu.scala 69:24]
  reg [31:0] DMemory_651; // @[cpu.scala 69:24]
  reg [31:0] DMemory_652; // @[cpu.scala 69:24]
  reg [31:0] DMemory_653; // @[cpu.scala 69:24]
  reg [31:0] DMemory_654; // @[cpu.scala 69:24]
  reg [31:0] DMemory_655; // @[cpu.scala 69:24]
  reg [31:0] DMemory_656; // @[cpu.scala 69:24]
  reg [31:0] DMemory_657; // @[cpu.scala 69:24]
  reg [31:0] DMemory_658; // @[cpu.scala 69:24]
  reg [31:0] DMemory_659; // @[cpu.scala 69:24]
  reg [31:0] DMemory_660; // @[cpu.scala 69:24]
  reg [31:0] DMemory_661; // @[cpu.scala 69:24]
  reg [31:0] DMemory_662; // @[cpu.scala 69:24]
  reg [31:0] DMemory_663; // @[cpu.scala 69:24]
  reg [31:0] DMemory_664; // @[cpu.scala 69:24]
  reg [31:0] DMemory_665; // @[cpu.scala 69:24]
  reg [31:0] DMemory_666; // @[cpu.scala 69:24]
  reg [31:0] DMemory_667; // @[cpu.scala 69:24]
  reg [31:0] DMemory_668; // @[cpu.scala 69:24]
  reg [31:0] DMemory_669; // @[cpu.scala 69:24]
  reg [31:0] DMemory_670; // @[cpu.scala 69:24]
  reg [31:0] DMemory_671; // @[cpu.scala 69:24]
  reg [31:0] DMemory_672; // @[cpu.scala 69:24]
  reg [31:0] DMemory_673; // @[cpu.scala 69:24]
  reg [31:0] DMemory_674; // @[cpu.scala 69:24]
  reg [31:0] DMemory_675; // @[cpu.scala 69:24]
  reg [31:0] DMemory_676; // @[cpu.scala 69:24]
  reg [31:0] DMemory_677; // @[cpu.scala 69:24]
  reg [31:0] DMemory_678; // @[cpu.scala 69:24]
  reg [31:0] DMemory_679; // @[cpu.scala 69:24]
  reg [31:0] DMemory_680; // @[cpu.scala 69:24]
  reg [31:0] DMemory_681; // @[cpu.scala 69:24]
  reg [31:0] DMemory_682; // @[cpu.scala 69:24]
  reg [31:0] DMemory_683; // @[cpu.scala 69:24]
  reg [31:0] DMemory_684; // @[cpu.scala 69:24]
  reg [31:0] DMemory_685; // @[cpu.scala 69:24]
  reg [31:0] DMemory_686; // @[cpu.scala 69:24]
  reg [31:0] DMemory_687; // @[cpu.scala 69:24]
  reg [31:0] DMemory_688; // @[cpu.scala 69:24]
  reg [31:0] DMemory_689; // @[cpu.scala 69:24]
  reg [31:0] DMemory_690; // @[cpu.scala 69:24]
  reg [31:0] DMemory_691; // @[cpu.scala 69:24]
  reg [31:0] DMemory_692; // @[cpu.scala 69:24]
  reg [31:0] DMemory_693; // @[cpu.scala 69:24]
  reg [31:0] DMemory_694; // @[cpu.scala 69:24]
  reg [31:0] DMemory_695; // @[cpu.scala 69:24]
  reg [31:0] DMemory_696; // @[cpu.scala 69:24]
  reg [31:0] DMemory_697; // @[cpu.scala 69:24]
  reg [31:0] DMemory_698; // @[cpu.scala 69:24]
  reg [31:0] DMemory_699; // @[cpu.scala 69:24]
  reg [31:0] DMemory_700; // @[cpu.scala 69:24]
  reg [31:0] DMemory_701; // @[cpu.scala 69:24]
  reg [31:0] DMemory_702; // @[cpu.scala 69:24]
  reg [31:0] DMemory_703; // @[cpu.scala 69:24]
  reg [31:0] DMemory_704; // @[cpu.scala 69:24]
  reg [31:0] DMemory_705; // @[cpu.scala 69:24]
  reg [31:0] DMemory_706; // @[cpu.scala 69:24]
  reg [31:0] DMemory_707; // @[cpu.scala 69:24]
  reg [31:0] DMemory_708; // @[cpu.scala 69:24]
  reg [31:0] DMemory_709; // @[cpu.scala 69:24]
  reg [31:0] DMemory_710; // @[cpu.scala 69:24]
  reg [31:0] DMemory_711; // @[cpu.scala 69:24]
  reg [31:0] DMemory_712; // @[cpu.scala 69:24]
  reg [31:0] DMemory_713; // @[cpu.scala 69:24]
  reg [31:0] DMemory_714; // @[cpu.scala 69:24]
  reg [31:0] DMemory_715; // @[cpu.scala 69:24]
  reg [31:0] DMemory_716; // @[cpu.scala 69:24]
  reg [31:0] DMemory_717; // @[cpu.scala 69:24]
  reg [31:0] DMemory_718; // @[cpu.scala 69:24]
  reg [31:0] DMemory_719; // @[cpu.scala 69:24]
  reg [31:0] DMemory_720; // @[cpu.scala 69:24]
  reg [31:0] DMemory_721; // @[cpu.scala 69:24]
  reg [31:0] DMemory_722; // @[cpu.scala 69:24]
  reg [31:0] DMemory_723; // @[cpu.scala 69:24]
  reg [31:0] DMemory_724; // @[cpu.scala 69:24]
  reg [31:0] DMemory_725; // @[cpu.scala 69:24]
  reg [31:0] DMemory_726; // @[cpu.scala 69:24]
  reg [31:0] DMemory_727; // @[cpu.scala 69:24]
  reg [31:0] DMemory_728; // @[cpu.scala 69:24]
  reg [31:0] DMemory_729; // @[cpu.scala 69:24]
  reg [31:0] DMemory_730; // @[cpu.scala 69:24]
  reg [31:0] DMemory_731; // @[cpu.scala 69:24]
  reg [31:0] DMemory_732; // @[cpu.scala 69:24]
  reg [31:0] DMemory_733; // @[cpu.scala 69:24]
  reg [31:0] DMemory_734; // @[cpu.scala 69:24]
  reg [31:0] DMemory_735; // @[cpu.scala 69:24]
  reg [31:0] DMemory_736; // @[cpu.scala 69:24]
  reg [31:0] DMemory_737; // @[cpu.scala 69:24]
  reg [31:0] DMemory_738; // @[cpu.scala 69:24]
  reg [31:0] DMemory_739; // @[cpu.scala 69:24]
  reg [31:0] DMemory_740; // @[cpu.scala 69:24]
  reg [31:0] DMemory_741; // @[cpu.scala 69:24]
  reg [31:0] DMemory_742; // @[cpu.scala 69:24]
  reg [31:0] DMemory_743; // @[cpu.scala 69:24]
  reg [31:0] DMemory_744; // @[cpu.scala 69:24]
  reg [31:0] DMemory_745; // @[cpu.scala 69:24]
  reg [31:0] DMemory_746; // @[cpu.scala 69:24]
  reg [31:0] DMemory_747; // @[cpu.scala 69:24]
  reg [31:0] DMemory_748; // @[cpu.scala 69:24]
  reg [31:0] DMemory_749; // @[cpu.scala 69:24]
  reg [31:0] DMemory_750; // @[cpu.scala 69:24]
  reg [31:0] DMemory_751; // @[cpu.scala 69:24]
  reg [31:0] DMemory_752; // @[cpu.scala 69:24]
  reg [31:0] DMemory_753; // @[cpu.scala 69:24]
  reg [31:0] DMemory_754; // @[cpu.scala 69:24]
  reg [31:0] DMemory_755; // @[cpu.scala 69:24]
  reg [31:0] DMemory_756; // @[cpu.scala 69:24]
  reg [31:0] DMemory_757; // @[cpu.scala 69:24]
  reg [31:0] DMemory_758; // @[cpu.scala 69:24]
  reg [31:0] DMemory_759; // @[cpu.scala 69:24]
  reg [31:0] DMemory_760; // @[cpu.scala 69:24]
  reg [31:0] DMemory_761; // @[cpu.scala 69:24]
  reg [31:0] DMemory_762; // @[cpu.scala 69:24]
  reg [31:0] DMemory_763; // @[cpu.scala 69:24]
  reg [31:0] DMemory_764; // @[cpu.scala 69:24]
  reg [31:0] DMemory_765; // @[cpu.scala 69:24]
  reg [31:0] DMemory_766; // @[cpu.scala 69:24]
  reg [31:0] DMemory_767; // @[cpu.scala 69:24]
  reg [31:0] DMemory_768; // @[cpu.scala 69:24]
  reg [31:0] DMemory_769; // @[cpu.scala 69:24]
  reg [31:0] DMemory_770; // @[cpu.scala 69:24]
  reg [31:0] DMemory_771; // @[cpu.scala 69:24]
  reg [31:0] DMemory_772; // @[cpu.scala 69:24]
  reg [31:0] DMemory_773; // @[cpu.scala 69:24]
  reg [31:0] DMemory_774; // @[cpu.scala 69:24]
  reg [31:0] DMemory_775; // @[cpu.scala 69:24]
  reg [31:0] DMemory_776; // @[cpu.scala 69:24]
  reg [31:0] DMemory_777; // @[cpu.scala 69:24]
  reg [31:0] DMemory_778; // @[cpu.scala 69:24]
  reg [31:0] DMemory_779; // @[cpu.scala 69:24]
  reg [31:0] DMemory_780; // @[cpu.scala 69:24]
  reg [31:0] DMemory_781; // @[cpu.scala 69:24]
  reg [31:0] DMemory_782; // @[cpu.scala 69:24]
  reg [31:0] DMemory_783; // @[cpu.scala 69:24]
  reg [31:0] DMemory_784; // @[cpu.scala 69:24]
  reg [31:0] DMemory_785; // @[cpu.scala 69:24]
  reg [31:0] DMemory_786; // @[cpu.scala 69:24]
  reg [31:0] DMemory_787; // @[cpu.scala 69:24]
  reg [31:0] DMemory_788; // @[cpu.scala 69:24]
  reg [31:0] DMemory_789; // @[cpu.scala 69:24]
  reg [31:0] DMemory_790; // @[cpu.scala 69:24]
  reg [31:0] DMemory_791; // @[cpu.scala 69:24]
  reg [31:0] DMemory_792; // @[cpu.scala 69:24]
  reg [31:0] DMemory_793; // @[cpu.scala 69:24]
  reg [31:0] DMemory_794; // @[cpu.scala 69:24]
  reg [31:0] DMemory_795; // @[cpu.scala 69:24]
  reg [31:0] DMemory_796; // @[cpu.scala 69:24]
  reg [31:0] DMemory_797; // @[cpu.scala 69:24]
  reg [31:0] DMemory_798; // @[cpu.scala 69:24]
  reg [31:0] DMemory_799; // @[cpu.scala 69:24]
  reg [31:0] DMemory_800; // @[cpu.scala 69:24]
  reg [31:0] DMemory_801; // @[cpu.scala 69:24]
  reg [31:0] DMemory_802; // @[cpu.scala 69:24]
  reg [31:0] DMemory_803; // @[cpu.scala 69:24]
  reg [31:0] DMemory_804; // @[cpu.scala 69:24]
  reg [31:0] DMemory_805; // @[cpu.scala 69:24]
  reg [31:0] DMemory_806; // @[cpu.scala 69:24]
  reg [31:0] DMemory_807; // @[cpu.scala 69:24]
  reg [31:0] DMemory_808; // @[cpu.scala 69:24]
  reg [31:0] DMemory_809; // @[cpu.scala 69:24]
  reg [31:0] DMemory_810; // @[cpu.scala 69:24]
  reg [31:0] DMemory_811; // @[cpu.scala 69:24]
  reg [31:0] DMemory_812; // @[cpu.scala 69:24]
  reg [31:0] DMemory_813; // @[cpu.scala 69:24]
  reg [31:0] DMemory_814; // @[cpu.scala 69:24]
  reg [31:0] DMemory_815; // @[cpu.scala 69:24]
  reg [31:0] DMemory_816; // @[cpu.scala 69:24]
  reg [31:0] DMemory_817; // @[cpu.scala 69:24]
  reg [31:0] DMemory_818; // @[cpu.scala 69:24]
  reg [31:0] DMemory_819; // @[cpu.scala 69:24]
  reg [31:0] DMemory_820; // @[cpu.scala 69:24]
  reg [31:0] DMemory_821; // @[cpu.scala 69:24]
  reg [31:0] DMemory_822; // @[cpu.scala 69:24]
  reg [31:0] DMemory_823; // @[cpu.scala 69:24]
  reg [31:0] DMemory_824; // @[cpu.scala 69:24]
  reg [31:0] DMemory_825; // @[cpu.scala 69:24]
  reg [31:0] DMemory_826; // @[cpu.scala 69:24]
  reg [31:0] DMemory_827; // @[cpu.scala 69:24]
  reg [31:0] DMemory_828; // @[cpu.scala 69:24]
  reg [31:0] DMemory_829; // @[cpu.scala 69:24]
  reg [31:0] DMemory_830; // @[cpu.scala 69:24]
  reg [31:0] DMemory_831; // @[cpu.scala 69:24]
  reg [31:0] DMemory_832; // @[cpu.scala 69:24]
  reg [31:0] DMemory_833; // @[cpu.scala 69:24]
  reg [31:0] DMemory_834; // @[cpu.scala 69:24]
  reg [31:0] DMemory_835; // @[cpu.scala 69:24]
  reg [31:0] DMemory_836; // @[cpu.scala 69:24]
  reg [31:0] DMemory_837; // @[cpu.scala 69:24]
  reg [31:0] DMemory_838; // @[cpu.scala 69:24]
  reg [31:0] DMemory_839; // @[cpu.scala 69:24]
  reg [31:0] DMemory_840; // @[cpu.scala 69:24]
  reg [31:0] DMemory_841; // @[cpu.scala 69:24]
  reg [31:0] DMemory_842; // @[cpu.scala 69:24]
  reg [31:0] DMemory_843; // @[cpu.scala 69:24]
  reg [31:0] DMemory_844; // @[cpu.scala 69:24]
  reg [31:0] DMemory_845; // @[cpu.scala 69:24]
  reg [31:0] DMemory_846; // @[cpu.scala 69:24]
  reg [31:0] DMemory_847; // @[cpu.scala 69:24]
  reg [31:0] DMemory_848; // @[cpu.scala 69:24]
  reg [31:0] DMemory_849; // @[cpu.scala 69:24]
  reg [31:0] DMemory_850; // @[cpu.scala 69:24]
  reg [31:0] DMemory_851; // @[cpu.scala 69:24]
  reg [31:0] DMemory_852; // @[cpu.scala 69:24]
  reg [31:0] DMemory_853; // @[cpu.scala 69:24]
  reg [31:0] DMemory_854; // @[cpu.scala 69:24]
  reg [31:0] DMemory_855; // @[cpu.scala 69:24]
  reg [31:0] DMemory_856; // @[cpu.scala 69:24]
  reg [31:0] DMemory_857; // @[cpu.scala 69:24]
  reg [31:0] DMemory_858; // @[cpu.scala 69:24]
  reg [31:0] DMemory_859; // @[cpu.scala 69:24]
  reg [31:0] DMemory_860; // @[cpu.scala 69:24]
  reg [31:0] DMemory_861; // @[cpu.scala 69:24]
  reg [31:0] DMemory_862; // @[cpu.scala 69:24]
  reg [31:0] DMemory_863; // @[cpu.scala 69:24]
  reg [31:0] DMemory_864; // @[cpu.scala 69:24]
  reg [31:0] DMemory_865; // @[cpu.scala 69:24]
  reg [31:0] DMemory_866; // @[cpu.scala 69:24]
  reg [31:0] DMemory_867; // @[cpu.scala 69:24]
  reg [31:0] DMemory_868; // @[cpu.scala 69:24]
  reg [31:0] DMemory_869; // @[cpu.scala 69:24]
  reg [31:0] DMemory_870; // @[cpu.scala 69:24]
  reg [31:0] DMemory_871; // @[cpu.scala 69:24]
  reg [31:0] DMemory_872; // @[cpu.scala 69:24]
  reg [31:0] DMemory_873; // @[cpu.scala 69:24]
  reg [31:0] DMemory_874; // @[cpu.scala 69:24]
  reg [31:0] DMemory_875; // @[cpu.scala 69:24]
  reg [31:0] DMemory_876; // @[cpu.scala 69:24]
  reg [31:0] DMemory_877; // @[cpu.scala 69:24]
  reg [31:0] DMemory_878; // @[cpu.scala 69:24]
  reg [31:0] DMemory_879; // @[cpu.scala 69:24]
  reg [31:0] DMemory_880; // @[cpu.scala 69:24]
  reg [31:0] DMemory_881; // @[cpu.scala 69:24]
  reg [31:0] DMemory_882; // @[cpu.scala 69:24]
  reg [31:0] DMemory_883; // @[cpu.scala 69:24]
  reg [31:0] DMemory_884; // @[cpu.scala 69:24]
  reg [31:0] DMemory_885; // @[cpu.scala 69:24]
  reg [31:0] DMemory_886; // @[cpu.scala 69:24]
  reg [31:0] DMemory_887; // @[cpu.scala 69:24]
  reg [31:0] DMemory_888; // @[cpu.scala 69:24]
  reg [31:0] DMemory_889; // @[cpu.scala 69:24]
  reg [31:0] DMemory_890; // @[cpu.scala 69:24]
  reg [31:0] DMemory_891; // @[cpu.scala 69:24]
  reg [31:0] DMemory_892; // @[cpu.scala 69:24]
  reg [31:0] DMemory_893; // @[cpu.scala 69:24]
  reg [31:0] DMemory_894; // @[cpu.scala 69:24]
  reg [31:0] DMemory_895; // @[cpu.scala 69:24]
  reg [31:0] DMemory_896; // @[cpu.scala 69:24]
  reg [31:0] DMemory_897; // @[cpu.scala 69:24]
  reg [31:0] DMemory_898; // @[cpu.scala 69:24]
  reg [31:0] DMemory_899; // @[cpu.scala 69:24]
  reg [31:0] DMemory_900; // @[cpu.scala 69:24]
  reg [31:0] DMemory_901; // @[cpu.scala 69:24]
  reg [31:0] DMemory_902; // @[cpu.scala 69:24]
  reg [31:0] DMemory_903; // @[cpu.scala 69:24]
  reg [31:0] DMemory_904; // @[cpu.scala 69:24]
  reg [31:0] DMemory_905; // @[cpu.scala 69:24]
  reg [31:0] DMemory_906; // @[cpu.scala 69:24]
  reg [31:0] DMemory_907; // @[cpu.scala 69:24]
  reg [31:0] DMemory_908; // @[cpu.scala 69:24]
  reg [31:0] DMemory_909; // @[cpu.scala 69:24]
  reg [31:0] DMemory_910; // @[cpu.scala 69:24]
  reg [31:0] DMemory_911; // @[cpu.scala 69:24]
  reg [31:0] DMemory_912; // @[cpu.scala 69:24]
  reg [31:0] DMemory_913; // @[cpu.scala 69:24]
  reg [31:0] DMemory_914; // @[cpu.scala 69:24]
  reg [31:0] DMemory_915; // @[cpu.scala 69:24]
  reg [31:0] DMemory_916; // @[cpu.scala 69:24]
  reg [31:0] DMemory_917; // @[cpu.scala 69:24]
  reg [31:0] DMemory_918; // @[cpu.scala 69:24]
  reg [31:0] DMemory_919; // @[cpu.scala 69:24]
  reg [31:0] DMemory_920; // @[cpu.scala 69:24]
  reg [31:0] DMemory_921; // @[cpu.scala 69:24]
  reg [31:0] DMemory_922; // @[cpu.scala 69:24]
  reg [31:0] DMemory_923; // @[cpu.scala 69:24]
  reg [31:0] DMemory_924; // @[cpu.scala 69:24]
  reg [31:0] DMemory_925; // @[cpu.scala 69:24]
  reg [31:0] DMemory_926; // @[cpu.scala 69:24]
  reg [31:0] DMemory_927; // @[cpu.scala 69:24]
  reg [31:0] DMemory_928; // @[cpu.scala 69:24]
  reg [31:0] DMemory_929; // @[cpu.scala 69:24]
  reg [31:0] DMemory_930; // @[cpu.scala 69:24]
  reg [31:0] DMemory_931; // @[cpu.scala 69:24]
  reg [31:0] DMemory_932; // @[cpu.scala 69:24]
  reg [31:0] DMemory_933; // @[cpu.scala 69:24]
  reg [31:0] DMemory_934; // @[cpu.scala 69:24]
  reg [31:0] DMemory_935; // @[cpu.scala 69:24]
  reg [31:0] DMemory_936; // @[cpu.scala 69:24]
  reg [31:0] DMemory_937; // @[cpu.scala 69:24]
  reg [31:0] DMemory_938; // @[cpu.scala 69:24]
  reg [31:0] DMemory_939; // @[cpu.scala 69:24]
  reg [31:0] DMemory_940; // @[cpu.scala 69:24]
  reg [31:0] DMemory_941; // @[cpu.scala 69:24]
  reg [31:0] DMemory_942; // @[cpu.scala 69:24]
  reg [31:0] DMemory_943; // @[cpu.scala 69:24]
  reg [31:0] DMemory_944; // @[cpu.scala 69:24]
  reg [31:0] DMemory_945; // @[cpu.scala 69:24]
  reg [31:0] DMemory_946; // @[cpu.scala 69:24]
  reg [31:0] DMemory_947; // @[cpu.scala 69:24]
  reg [31:0] DMemory_948; // @[cpu.scala 69:24]
  reg [31:0] DMemory_949; // @[cpu.scala 69:24]
  reg [31:0] DMemory_950; // @[cpu.scala 69:24]
  reg [31:0] DMemory_951; // @[cpu.scala 69:24]
  reg [31:0] DMemory_952; // @[cpu.scala 69:24]
  reg [31:0] DMemory_953; // @[cpu.scala 69:24]
  reg [31:0] DMemory_954; // @[cpu.scala 69:24]
  reg [31:0] DMemory_955; // @[cpu.scala 69:24]
  reg [31:0] DMemory_956; // @[cpu.scala 69:24]
  reg [31:0] DMemory_957; // @[cpu.scala 69:24]
  reg [31:0] DMemory_958; // @[cpu.scala 69:24]
  reg [31:0] DMemory_959; // @[cpu.scala 69:24]
  reg [31:0] DMemory_960; // @[cpu.scala 69:24]
  reg [31:0] DMemory_961; // @[cpu.scala 69:24]
  reg [31:0] DMemory_962; // @[cpu.scala 69:24]
  reg [31:0] DMemory_963; // @[cpu.scala 69:24]
  reg [31:0] DMemory_964; // @[cpu.scala 69:24]
  reg [31:0] DMemory_965; // @[cpu.scala 69:24]
  reg [31:0] DMemory_966; // @[cpu.scala 69:24]
  reg [31:0] DMemory_967; // @[cpu.scala 69:24]
  reg [31:0] DMemory_968; // @[cpu.scala 69:24]
  reg [31:0] DMemory_969; // @[cpu.scala 69:24]
  reg [31:0] DMemory_970; // @[cpu.scala 69:24]
  reg [31:0] DMemory_971; // @[cpu.scala 69:24]
  reg [31:0] DMemory_972; // @[cpu.scala 69:24]
  reg [31:0] DMemory_973; // @[cpu.scala 69:24]
  reg [31:0] DMemory_974; // @[cpu.scala 69:24]
  reg [31:0] DMemory_975; // @[cpu.scala 69:24]
  reg [31:0] DMemory_976; // @[cpu.scala 69:24]
  reg [31:0] DMemory_977; // @[cpu.scala 69:24]
  reg [31:0] DMemory_978; // @[cpu.scala 69:24]
  reg [31:0] DMemory_979; // @[cpu.scala 69:24]
  reg [31:0] DMemory_980; // @[cpu.scala 69:24]
  reg [31:0] DMemory_981; // @[cpu.scala 69:24]
  reg [31:0] DMemory_982; // @[cpu.scala 69:24]
  reg [31:0] DMemory_983; // @[cpu.scala 69:24]
  reg [31:0] DMemory_984; // @[cpu.scala 69:24]
  reg [31:0] DMemory_985; // @[cpu.scala 69:24]
  reg [31:0] DMemory_986; // @[cpu.scala 69:24]
  reg [31:0] DMemory_987; // @[cpu.scala 69:24]
  reg [31:0] DMemory_988; // @[cpu.scala 69:24]
  reg [31:0] DMemory_989; // @[cpu.scala 69:24]
  reg [31:0] DMemory_990; // @[cpu.scala 69:24]
  reg [31:0] DMemory_991; // @[cpu.scala 69:24]
  reg [31:0] DMemory_992; // @[cpu.scala 69:24]
  reg [31:0] DMemory_993; // @[cpu.scala 69:24]
  reg [31:0] DMemory_994; // @[cpu.scala 69:24]
  reg [31:0] DMemory_995; // @[cpu.scala 69:24]
  reg [31:0] DMemory_996; // @[cpu.scala 69:24]
  reg [31:0] DMemory_997; // @[cpu.scala 69:24]
  reg [31:0] DMemory_998; // @[cpu.scala 69:24]
  reg [31:0] DMemory_999; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1000; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1001; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1002; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1003; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1004; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1005; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1006; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1007; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1008; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1009; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1010; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1011; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1012; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1013; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1014; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1015; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1016; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1017; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1018; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1019; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1020; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1021; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1022; // @[cpu.scala 69:24]
  reg [31:0] DMemory_1023; // @[cpu.scala 69:24]
  reg [31:0] IMemory_0; // @[cpu.scala 70:24]
  reg [31:0] IMemory_1; // @[cpu.scala 70:24]
  reg [31:0] IFIDIR; // @[cpu.scala 73:49]
  reg [31:0] IDEXIR; // @[cpu.scala 73:49]
  reg [31:0] EXMEMIR; // @[cpu.scala 73:49]
  reg [31:0] MEMWBIR; // @[cpu.scala 73:49]
  reg [63:0] CurPC; // @[cpu.scala 76:22]
  wire [4:0] EXMEMrd = EXMEMIR[11:7]; // @[cpu.scala 105:32]
  wire [4:0] IDEXrd = IDEXIR[11:7]; // @[cpu.scala 106:30]
  wire [2:0] IFID_funct3 = IFIDIR[14:12]; // @[cpu.scala 107:29]
  wire [4:0] IFIDrs1 = io_rvfi_rst ? IFIDIR[19:15] : IFIDIR[19:15]; // @[cpu.scala 80:21 82:13 97:13]
  wire [4:0] MEMWBrd = io_rvfi_rst ? MEMWBIR[11:7] : MEMWBIR[11:7]; // @[cpu.scala 103:13 80:21 88:13]
  wire  _bypassAFromWB_T_1 = IFIDrs1 != 5'h0; // @[cpu.scala 110:41]
  wire [6:0] MEMWBop = io_rvfi_rst ? MEMWBIR[6:0] : MEMWBIR[6:0]; // @[cpu.scala 102:13 80:21 87:13]
  wire  _bypassAFromWB_T_3 = MEMWBop == 7'h33; // @[cpu.scala 110:62]
  wire  _bypassAFromWB_T_4 = MEMWBop == 7'h3; // @[cpu.scala 110:83]
  wire  _bypassAFromWB_T_5 = MEMWBop == 7'h33 | MEMWBop == 7'h3; // @[cpu.scala 110:72]
  wire  bypassAFromWB = IFIDrs1 == MEMWBrd & IFIDrs1 != 5'h0 & (MEMWBop == 7'h33 | MEMWBop == 7'h3); // @[cpu.scala 110:50]
  wire [4:0] IFIDrs2 = io_rvfi_rst ? IFIDIR[24:20] : IFIDIR[24:20]; // @[cpu.scala 80:21 83:13 98:13]
  wire  _bypassBFromWB_T_1 = IFIDrs2 != 5'h0; // @[cpu.scala 112:41]
  wire  bypassBFromWB = IFIDrs2 == MEMWBrd & IFIDrs2 != 5'h0 & _bypassAFromWB_T_5; // @[cpu.scala 112:50]
  wire  _bypassAFromMEM_T_2 = IFIDrs1 == EXMEMrd & _bypassAFromWB_T_1; // @[cpu.scala 114:29]
  wire [6:0] EXMEMop = io_rvfi_rst ? EXMEMIR[6:0] : EXMEMIR[6:0]; // @[cpu.scala 101:13 80:21 86:13]
  wire  _bypassAFromMEM_T_3 = EXMEMop == 7'h33; // @[cpu.scala 114:62]
  wire  bypassAFromMEM = IFIDrs1 == EXMEMrd & _bypassAFromWB_T_1 & EXMEMop == 7'h33; // @[cpu.scala 114:50]
  wire  _bypassBFromMEM_T_2 = IFIDrs2 == EXMEMrd & _bypassBFromWB_T_1; // @[cpu.scala 116:29]
  wire  bypassBFromMEM = IFIDrs2 == EXMEMrd & _bypassBFromWB_T_1 & _bypassAFromMEM_T_3; // @[cpu.scala 116:50]
  wire  _bypassAFromEX_T_2 = IFIDrs1 == IDEXrd & _bypassAFromWB_T_1; // @[cpu.scala 118:28]
  wire [6:0] IDEXop = io_rvfi_rst ? IDEXIR[6:0] : IDEXIR[6:0]; // @[cpu.scala 80:21 84:12 99:12]
  wire  _bypassAFromEX_T_3 = IDEXop == 7'h33; // @[cpu.scala 118:60]
  wire  bypassAFromEX = IFIDrs1 == IDEXrd & _bypassAFromWB_T_1 & IDEXop == 7'h33; // @[cpu.scala 118:49]
  wire  _bypassBFromEX_T_2 = IFIDrs2 == IDEXrd & _bypassBFromWB_T_1; // @[cpu.scala 120:28]
  wire  bypassBFromEX = IFIDrs2 == IDEXrd & _bypassBFromWB_T_1 & _bypassAFromEX_T_3; // @[cpu.scala 120:49]
  wire  _stall_T = EXMEMop == 7'h3; // @[cpu.scala 123:16]
  wire  _stall_T_8 = EXMEMop == 7'h3 & (_bypassAFromMEM_T_2 | _bypassBFromMEM_T_2); // @[cpu.scala 123:24]
  wire  _stall_T_9 = IDEXop == 7'h3; // @[cpu.scala 125:15]
  wire  _stall_T_17 = IDEXop == 7'h3 & (_bypassAFromEX_T_2 | _bypassBFromEX_T_2); // @[cpu.scala 125:23]
  wire  stall = _stall_T_8 | _stall_T_17; // @[cpu.scala 124:7]
  wire [6:0] IFIDop = io_rvfi_rst ? IFIDIR[6:0] : IFIDIR[6:0]; // @[cpu.scala 100:12 80:21 85:12]
  wire [63:0] _A_T_1 = IDEXA + IDEXB; // @[cpu.scala 166:20]
  wire [63:0] _GEN_1029 = 5'h1 == IFIDrs1 ? Regs_1 : Regs_0; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1030 = 5'h2 == IFIDrs1 ? Regs_2 : _GEN_1029; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1031 = 5'h3 == IFIDrs1 ? Regs_3 : _GEN_1030; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1032 = 5'h4 == IFIDrs1 ? Regs_4 : _GEN_1031; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1033 = 5'h5 == IFIDrs1 ? Regs_5 : _GEN_1032; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1034 = 5'h6 == IFIDrs1 ? Regs_6 : _GEN_1033; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1035 = 5'h7 == IFIDrs1 ? Regs_7 : _GEN_1034; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1036 = 5'h8 == IFIDrs1 ? Regs_8 : _GEN_1035; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1037 = 5'h9 == IFIDrs1 ? Regs_9 : _GEN_1036; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1038 = 5'ha == IFIDrs1 ? Regs_10 : _GEN_1037; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1039 = 5'hb == IFIDrs1 ? Regs_11 : _GEN_1038; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1040 = 5'hc == IFIDrs1 ? Regs_12 : _GEN_1039; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1041 = 5'hd == IFIDrs1 ? Regs_13 : _GEN_1040; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1042 = 5'he == IFIDrs1 ? Regs_14 : _GEN_1041; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1043 = 5'hf == IFIDrs1 ? Regs_15 : _GEN_1042; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1044 = 5'h10 == IFIDrs1 ? Regs_16 : _GEN_1043; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1045 = 5'h11 == IFIDrs1 ? Regs_17 : _GEN_1044; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1046 = 5'h12 == IFIDrs1 ? Regs_18 : _GEN_1045; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1047 = 5'h13 == IFIDrs1 ? Regs_19 : _GEN_1046; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1048 = 5'h14 == IFIDrs1 ? Regs_20 : _GEN_1047; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1049 = 5'h15 == IFIDrs1 ? Regs_21 : _GEN_1048; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1050 = 5'h16 == IFIDrs1 ? Regs_22 : _GEN_1049; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1051 = 5'h17 == IFIDrs1 ? Regs_23 : _GEN_1050; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1052 = 5'h18 == IFIDrs1 ? Regs_24 : _GEN_1051; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1053 = 5'h19 == IFIDrs1 ? Regs_25 : _GEN_1052; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1054 = 5'h1a == IFIDrs1 ? Regs_26 : _GEN_1053; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1055 = 5'h1b == IFIDrs1 ? Regs_27 : _GEN_1054; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1056 = 5'h1c == IFIDrs1 ? Regs_28 : _GEN_1055; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1057 = 5'h1d == IFIDrs1 ? Regs_29 : _GEN_1056; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1058 = 5'h1e == IFIDrs1 ? Regs_30 : _GEN_1057; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1059 = 5'h1f == IFIDrs1 ? Regs_31 : _GEN_1058; // @[cpu.scala 174:{15,15}]
  wire [63:0] _GEN_1061 = bypassAFromWB ? MEMWBValue : _GEN_1059; // @[cpu.scala 170:33 172:11 175:11]
  wire [63:0] _GEN_1063 = bypassAFromMEM ? EXMEMALUOut : _GEN_1061; // @[cpu.scala 167:34 169:11]
  wire [63:0] _GEN_1065 = bypassAFromEX ? _A_T_1 : _GEN_1063; // @[cpu.scala 164:27 166:11]
  wire [63:0] A = ~stall ? _GEN_1065 : 64'h0; // @[cpu.scala 137:27]
  wire [63:0] _B_T_1 = IDEXB + IDEXA; // @[cpu.scala 179:20]
  wire [63:0] _GEN_1067 = 5'h1 == IFIDrs2 ? Regs_1 : Regs_0; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1068 = 5'h2 == IFIDrs2 ? Regs_2 : _GEN_1067; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1069 = 5'h3 == IFIDrs2 ? Regs_3 : _GEN_1068; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1070 = 5'h4 == IFIDrs2 ? Regs_4 : _GEN_1069; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1071 = 5'h5 == IFIDrs2 ? Regs_5 : _GEN_1070; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1072 = 5'h6 == IFIDrs2 ? Regs_6 : _GEN_1071; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1073 = 5'h7 == IFIDrs2 ? Regs_7 : _GEN_1072; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1074 = 5'h8 == IFIDrs2 ? Regs_8 : _GEN_1073; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1075 = 5'h9 == IFIDrs2 ? Regs_9 : _GEN_1074; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1076 = 5'ha == IFIDrs2 ? Regs_10 : _GEN_1075; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1077 = 5'hb == IFIDrs2 ? Regs_11 : _GEN_1076; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1078 = 5'hc == IFIDrs2 ? Regs_12 : _GEN_1077; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1079 = 5'hd == IFIDrs2 ? Regs_13 : _GEN_1078; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1080 = 5'he == IFIDrs2 ? Regs_14 : _GEN_1079; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1081 = 5'hf == IFIDrs2 ? Regs_15 : _GEN_1080; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1082 = 5'h10 == IFIDrs2 ? Regs_16 : _GEN_1081; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1083 = 5'h11 == IFIDrs2 ? Regs_17 : _GEN_1082; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1084 = 5'h12 == IFIDrs2 ? Regs_18 : _GEN_1083; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1085 = 5'h13 == IFIDrs2 ? Regs_19 : _GEN_1084; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1086 = 5'h14 == IFIDrs2 ? Regs_20 : _GEN_1085; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1087 = 5'h15 == IFIDrs2 ? Regs_21 : _GEN_1086; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1088 = 5'h16 == IFIDrs2 ? Regs_22 : _GEN_1087; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1089 = 5'h17 == IFIDrs2 ? Regs_23 : _GEN_1088; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1090 = 5'h18 == IFIDrs2 ? Regs_24 : _GEN_1089; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1091 = 5'h19 == IFIDrs2 ? Regs_25 : _GEN_1090; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1092 = 5'h1a == IFIDrs2 ? Regs_26 : _GEN_1091; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1093 = 5'h1b == IFIDrs2 ? Regs_27 : _GEN_1092; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1094 = 5'h1c == IFIDrs2 ? Regs_28 : _GEN_1093; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1095 = 5'h1d == IFIDrs2 ? Regs_29 : _GEN_1094; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1096 = 5'h1e == IFIDrs2 ? Regs_30 : _GEN_1095; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1097 = 5'h1f == IFIDrs2 ? Regs_31 : _GEN_1096; // @[cpu.scala 187:{15,15}]
  wire [63:0] _GEN_1099 = bypassBFromWB ? MEMWBValue : _GEN_1097; // @[cpu.scala 183:33 185:11 188:11]
  wire [63:0] _GEN_1101 = bypassBFromMEM ? EXMEMALUOut : _GEN_1099; // @[cpu.scala 180:34 182:11]
  wire [63:0] _GEN_1103 = bypassBFromEX ? _B_T_1 : _GEN_1101; // @[cpu.scala 177:27 179:11]
  wire [63:0] B = ~stall ? _GEN_1103 : 64'h0; // @[cpu.scala 137:27]
  wire  takeBranch = IFIDop == 7'h63 & IFID_funct3 == 3'h0 & A == B; // @[cpu.scala 129:64]
  wire [63:0] _IFIDIR_T = {{2'd0}, PC[63:2]}; // @[cpu.scala 141:31]
  wire [31:0] _GEN_1 = 10'h1 == _IFIDIR_T[9:0] ? IMemory_1 : IMemory_0; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_2 = 10'h2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_3 = 10'h3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_2; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_4 = 10'h4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_3; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_5 = 10'h5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_4; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_6 = 10'h6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_5; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_7 = 10'h7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_6; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_8 = 10'h8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_7; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_9 = 10'h9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_8; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_10 = 10'ha == _IFIDIR_T[9:0] ? 32'h13 : _GEN_9; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_11 = 10'hb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_10; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_12 = 10'hc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_11; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_13 = 10'hd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_12; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_14 = 10'he == _IFIDIR_T[9:0] ? 32'h13 : _GEN_13; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_15 = 10'hf == _IFIDIR_T[9:0] ? 32'h13 : _GEN_14; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_16 = 10'h10 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_15; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_17 = 10'h11 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_16; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_18 = 10'h12 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_17; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_19 = 10'h13 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_18; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_20 = 10'h14 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_19; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_21 = 10'h15 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_20; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_22 = 10'h16 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_21; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_23 = 10'h17 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_22; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_24 = 10'h18 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_23; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_25 = 10'h19 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_24; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_26 = 10'h1a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_25; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_27 = 10'h1b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_26; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_28 = 10'h1c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_27; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_29 = 10'h1d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_28; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_30 = 10'h1e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_29; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_31 = 10'h1f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_30; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_32 = 10'h20 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_31; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_33 = 10'h21 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_32; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_34 = 10'h22 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_33; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_35 = 10'h23 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_34; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_36 = 10'h24 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_35; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_37 = 10'h25 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_36; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_38 = 10'h26 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_37; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_39 = 10'h27 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_38; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_40 = 10'h28 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_39; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_41 = 10'h29 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_40; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_42 = 10'h2a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_41; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_43 = 10'h2b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_42; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_44 = 10'h2c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_43; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_45 = 10'h2d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_44; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_46 = 10'h2e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_45; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_47 = 10'h2f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_46; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_48 = 10'h30 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_47; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_49 = 10'h31 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_48; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_50 = 10'h32 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_49; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_51 = 10'h33 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_50; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_52 = 10'h34 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_51; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_53 = 10'h35 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_52; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_54 = 10'h36 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_53; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_55 = 10'h37 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_54; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_56 = 10'h38 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_55; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_57 = 10'h39 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_56; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_58 = 10'h3a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_57; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_59 = 10'h3b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_58; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_60 = 10'h3c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_59; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_61 = 10'h3d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_60; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_62 = 10'h3e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_61; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_63 = 10'h3f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_62; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_64 = 10'h40 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_63; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_65 = 10'h41 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_64; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_66 = 10'h42 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_65; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_67 = 10'h43 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_66; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_68 = 10'h44 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_67; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_69 = 10'h45 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_68; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_70 = 10'h46 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_69; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_71 = 10'h47 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_70; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_72 = 10'h48 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_71; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_73 = 10'h49 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_72; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_74 = 10'h4a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_73; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_75 = 10'h4b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_74; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_76 = 10'h4c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_75; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_77 = 10'h4d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_76; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_78 = 10'h4e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_77; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_79 = 10'h4f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_78; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_80 = 10'h50 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_79; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_81 = 10'h51 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_80; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_82 = 10'h52 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_81; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_83 = 10'h53 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_82; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_84 = 10'h54 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_83; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_85 = 10'h55 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_84; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_86 = 10'h56 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_85; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_87 = 10'h57 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_86; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_88 = 10'h58 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_87; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_89 = 10'h59 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_88; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_90 = 10'h5a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_89; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_91 = 10'h5b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_90; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_92 = 10'h5c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_91; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_93 = 10'h5d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_92; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_94 = 10'h5e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_93; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_95 = 10'h5f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_94; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_96 = 10'h60 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_95; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_97 = 10'h61 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_96; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_98 = 10'h62 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_97; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_99 = 10'h63 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_98; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_100 = 10'h64 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_99; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_101 = 10'h65 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_100; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_102 = 10'h66 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_101; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_103 = 10'h67 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_102; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_104 = 10'h68 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_103; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_105 = 10'h69 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_104; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_106 = 10'h6a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_105; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_107 = 10'h6b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_106; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_108 = 10'h6c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_107; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_109 = 10'h6d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_108; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_110 = 10'h6e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_109; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_111 = 10'h6f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_110; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_112 = 10'h70 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_111; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_113 = 10'h71 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_112; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_114 = 10'h72 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_113; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_115 = 10'h73 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_114; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_116 = 10'h74 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_115; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_117 = 10'h75 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_116; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_118 = 10'h76 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_117; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_119 = 10'h77 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_118; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_120 = 10'h78 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_119; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_121 = 10'h79 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_120; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_122 = 10'h7a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_121; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_123 = 10'h7b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_122; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_124 = 10'h7c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_123; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_125 = 10'h7d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_124; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_126 = 10'h7e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_125; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_127 = 10'h7f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_126; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_128 = 10'h80 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_127; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_129 = 10'h81 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_128; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_130 = 10'h82 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_129; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_131 = 10'h83 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_130; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_132 = 10'h84 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_131; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_133 = 10'h85 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_132; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_134 = 10'h86 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_133; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_135 = 10'h87 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_134; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_136 = 10'h88 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_135; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_137 = 10'h89 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_136; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_138 = 10'h8a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_137; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_139 = 10'h8b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_138; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_140 = 10'h8c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_139; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_141 = 10'h8d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_140; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_142 = 10'h8e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_141; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_143 = 10'h8f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_142; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_144 = 10'h90 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_143; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_145 = 10'h91 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_144; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_146 = 10'h92 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_145; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_147 = 10'h93 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_146; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_148 = 10'h94 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_147; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_149 = 10'h95 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_148; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_150 = 10'h96 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_149; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_151 = 10'h97 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_150; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_152 = 10'h98 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_151; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_153 = 10'h99 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_152; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_154 = 10'h9a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_153; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_155 = 10'h9b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_154; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_156 = 10'h9c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_155; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_157 = 10'h9d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_156; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_158 = 10'h9e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_157; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_159 = 10'h9f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_158; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_160 = 10'ha0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_159; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_161 = 10'ha1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_160; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_162 = 10'ha2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_161; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_163 = 10'ha3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_162; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_164 = 10'ha4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_163; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_165 = 10'ha5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_164; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_166 = 10'ha6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_165; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_167 = 10'ha7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_166; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_168 = 10'ha8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_167; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_169 = 10'ha9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_168; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_170 = 10'haa == _IFIDIR_T[9:0] ? 32'h13 : _GEN_169; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_171 = 10'hab == _IFIDIR_T[9:0] ? 32'h13 : _GEN_170; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_172 = 10'hac == _IFIDIR_T[9:0] ? 32'h13 : _GEN_171; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_173 = 10'had == _IFIDIR_T[9:0] ? 32'h13 : _GEN_172; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_174 = 10'hae == _IFIDIR_T[9:0] ? 32'h13 : _GEN_173; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_175 = 10'haf == _IFIDIR_T[9:0] ? 32'h13 : _GEN_174; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_176 = 10'hb0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_175; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_177 = 10'hb1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_176; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_178 = 10'hb2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_177; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_179 = 10'hb3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_178; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_180 = 10'hb4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_179; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_181 = 10'hb5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_180; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_182 = 10'hb6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_181; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_183 = 10'hb7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_182; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_184 = 10'hb8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_183; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_185 = 10'hb9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_184; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_186 = 10'hba == _IFIDIR_T[9:0] ? 32'h13 : _GEN_185; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_187 = 10'hbb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_186; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_188 = 10'hbc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_187; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_189 = 10'hbd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_188; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_190 = 10'hbe == _IFIDIR_T[9:0] ? 32'h13 : _GEN_189; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_191 = 10'hbf == _IFIDIR_T[9:0] ? 32'h13 : _GEN_190; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_192 = 10'hc0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_191; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_193 = 10'hc1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_192; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_194 = 10'hc2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_193; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_195 = 10'hc3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_194; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_196 = 10'hc4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_195; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_197 = 10'hc5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_196; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_198 = 10'hc6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_197; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_199 = 10'hc7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_198; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_200 = 10'hc8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_199; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_201 = 10'hc9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_200; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_202 = 10'hca == _IFIDIR_T[9:0] ? 32'h13 : _GEN_201; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_203 = 10'hcb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_202; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_204 = 10'hcc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_203; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_205 = 10'hcd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_204; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_206 = 10'hce == _IFIDIR_T[9:0] ? 32'h13 : _GEN_205; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_207 = 10'hcf == _IFIDIR_T[9:0] ? 32'h13 : _GEN_206; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_208 = 10'hd0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_207; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_209 = 10'hd1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_208; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_210 = 10'hd2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_209; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_211 = 10'hd3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_210; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_212 = 10'hd4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_211; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_213 = 10'hd5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_212; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_214 = 10'hd6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_213; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_215 = 10'hd7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_214; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_216 = 10'hd8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_215; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_217 = 10'hd9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_216; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_218 = 10'hda == _IFIDIR_T[9:0] ? 32'h13 : _GEN_217; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_219 = 10'hdb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_218; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_220 = 10'hdc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_219; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_221 = 10'hdd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_220; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_222 = 10'hde == _IFIDIR_T[9:0] ? 32'h13 : _GEN_221; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_223 = 10'hdf == _IFIDIR_T[9:0] ? 32'h13 : _GEN_222; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_224 = 10'he0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_223; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_225 = 10'he1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_224; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_226 = 10'he2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_225; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_227 = 10'he3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_226; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_228 = 10'he4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_227; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_229 = 10'he5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_228; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_230 = 10'he6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_229; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_231 = 10'he7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_230; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_232 = 10'he8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_231; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_233 = 10'he9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_232; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_234 = 10'hea == _IFIDIR_T[9:0] ? 32'h13 : _GEN_233; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_235 = 10'heb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_234; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_236 = 10'hec == _IFIDIR_T[9:0] ? 32'h13 : _GEN_235; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_237 = 10'hed == _IFIDIR_T[9:0] ? 32'h13 : _GEN_236; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_238 = 10'hee == _IFIDIR_T[9:0] ? 32'h13 : _GEN_237; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_239 = 10'hef == _IFIDIR_T[9:0] ? 32'h13 : _GEN_238; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_240 = 10'hf0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_239; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_241 = 10'hf1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_240; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_242 = 10'hf2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_241; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_243 = 10'hf3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_242; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_244 = 10'hf4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_243; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_245 = 10'hf5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_244; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_246 = 10'hf6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_245; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_247 = 10'hf7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_246; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_248 = 10'hf8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_247; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_249 = 10'hf9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_248; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_250 = 10'hfa == _IFIDIR_T[9:0] ? 32'h13 : _GEN_249; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_251 = 10'hfb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_250; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_252 = 10'hfc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_251; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_253 = 10'hfd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_252; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_254 = 10'hfe == _IFIDIR_T[9:0] ? 32'h13 : _GEN_253; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_255 = 10'hff == _IFIDIR_T[9:0] ? 32'h13 : _GEN_254; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_256 = 10'h100 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_255; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_257 = 10'h101 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_256; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_258 = 10'h102 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_257; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_259 = 10'h103 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_258; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_260 = 10'h104 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_259; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_261 = 10'h105 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_260; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_262 = 10'h106 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_261; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_263 = 10'h107 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_262; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_264 = 10'h108 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_263; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_265 = 10'h109 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_264; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_266 = 10'h10a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_265; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_267 = 10'h10b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_266; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_268 = 10'h10c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_267; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_269 = 10'h10d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_268; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_270 = 10'h10e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_269; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_271 = 10'h10f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_270; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_272 = 10'h110 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_271; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_273 = 10'h111 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_272; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_274 = 10'h112 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_273; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_275 = 10'h113 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_274; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_276 = 10'h114 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_275; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_277 = 10'h115 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_276; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_278 = 10'h116 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_277; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_279 = 10'h117 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_278; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_280 = 10'h118 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_279; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_281 = 10'h119 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_280; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_282 = 10'h11a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_281; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_283 = 10'h11b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_282; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_284 = 10'h11c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_283; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_285 = 10'h11d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_284; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_286 = 10'h11e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_285; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_287 = 10'h11f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_286; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_288 = 10'h120 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_287; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_289 = 10'h121 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_288; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_290 = 10'h122 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_289; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_291 = 10'h123 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_290; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_292 = 10'h124 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_291; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_293 = 10'h125 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_292; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_294 = 10'h126 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_293; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_295 = 10'h127 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_294; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_296 = 10'h128 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_295; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_297 = 10'h129 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_296; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_298 = 10'h12a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_297; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_299 = 10'h12b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_298; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_300 = 10'h12c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_299; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_301 = 10'h12d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_300; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_302 = 10'h12e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_301; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_303 = 10'h12f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_302; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_304 = 10'h130 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_303; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_305 = 10'h131 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_304; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_306 = 10'h132 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_305; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_307 = 10'h133 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_306; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_308 = 10'h134 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_307; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_309 = 10'h135 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_308; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_310 = 10'h136 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_309; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_311 = 10'h137 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_310; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_312 = 10'h138 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_311; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_313 = 10'h139 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_312; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_314 = 10'h13a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_313; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_315 = 10'h13b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_314; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_316 = 10'h13c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_315; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_317 = 10'h13d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_316; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_318 = 10'h13e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_317; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_319 = 10'h13f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_318; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_320 = 10'h140 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_319; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_321 = 10'h141 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_320; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_322 = 10'h142 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_321; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_323 = 10'h143 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_322; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_324 = 10'h144 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_323; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_325 = 10'h145 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_324; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_326 = 10'h146 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_325; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_327 = 10'h147 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_326; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_328 = 10'h148 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_327; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_329 = 10'h149 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_328; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_330 = 10'h14a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_329; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_331 = 10'h14b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_330; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_332 = 10'h14c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_331; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_333 = 10'h14d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_332; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_334 = 10'h14e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_333; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_335 = 10'h14f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_334; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_336 = 10'h150 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_335; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_337 = 10'h151 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_336; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_338 = 10'h152 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_337; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_339 = 10'h153 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_338; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_340 = 10'h154 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_339; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_341 = 10'h155 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_340; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_342 = 10'h156 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_341; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_343 = 10'h157 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_342; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_344 = 10'h158 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_343; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_345 = 10'h159 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_344; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_346 = 10'h15a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_345; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_347 = 10'h15b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_346; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_348 = 10'h15c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_347; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_349 = 10'h15d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_348; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_350 = 10'h15e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_349; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_351 = 10'h15f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_350; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_352 = 10'h160 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_351; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_353 = 10'h161 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_352; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_354 = 10'h162 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_353; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_355 = 10'h163 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_354; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_356 = 10'h164 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_355; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_357 = 10'h165 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_356; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_358 = 10'h166 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_357; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_359 = 10'h167 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_358; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_360 = 10'h168 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_359; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_361 = 10'h169 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_360; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_362 = 10'h16a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_361; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_363 = 10'h16b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_362; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_364 = 10'h16c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_363; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_365 = 10'h16d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_364; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_366 = 10'h16e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_365; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_367 = 10'h16f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_366; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_368 = 10'h170 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_367; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_369 = 10'h171 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_368; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_370 = 10'h172 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_369; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_371 = 10'h173 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_370; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_372 = 10'h174 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_371; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_373 = 10'h175 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_372; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_374 = 10'h176 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_373; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_375 = 10'h177 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_374; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_376 = 10'h178 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_375; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_377 = 10'h179 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_376; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_378 = 10'h17a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_377; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_379 = 10'h17b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_378; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_380 = 10'h17c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_379; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_381 = 10'h17d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_380; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_382 = 10'h17e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_381; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_383 = 10'h17f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_382; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_384 = 10'h180 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_383; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_385 = 10'h181 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_384; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_386 = 10'h182 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_385; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_387 = 10'h183 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_386; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_388 = 10'h184 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_387; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_389 = 10'h185 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_388; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_390 = 10'h186 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_389; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_391 = 10'h187 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_390; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_392 = 10'h188 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_391; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_393 = 10'h189 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_392; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_394 = 10'h18a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_393; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_395 = 10'h18b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_394; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_396 = 10'h18c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_395; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_397 = 10'h18d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_396; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_398 = 10'h18e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_397; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_399 = 10'h18f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_398; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_400 = 10'h190 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_399; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_401 = 10'h191 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_400; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_402 = 10'h192 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_401; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_403 = 10'h193 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_402; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_404 = 10'h194 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_403; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_405 = 10'h195 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_404; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_406 = 10'h196 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_405; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_407 = 10'h197 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_406; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_408 = 10'h198 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_407; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_409 = 10'h199 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_408; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_410 = 10'h19a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_409; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_411 = 10'h19b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_410; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_412 = 10'h19c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_411; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_413 = 10'h19d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_412; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_414 = 10'h19e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_413; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_415 = 10'h19f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_414; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_416 = 10'h1a0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_415; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_417 = 10'h1a1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_416; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_418 = 10'h1a2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_417; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_419 = 10'h1a3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_418; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_420 = 10'h1a4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_419; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_421 = 10'h1a5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_420; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_422 = 10'h1a6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_421; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_423 = 10'h1a7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_422; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_424 = 10'h1a8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_423; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_425 = 10'h1a9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_424; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_426 = 10'h1aa == _IFIDIR_T[9:0] ? 32'h13 : _GEN_425; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_427 = 10'h1ab == _IFIDIR_T[9:0] ? 32'h13 : _GEN_426; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_428 = 10'h1ac == _IFIDIR_T[9:0] ? 32'h13 : _GEN_427; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_429 = 10'h1ad == _IFIDIR_T[9:0] ? 32'h13 : _GEN_428; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_430 = 10'h1ae == _IFIDIR_T[9:0] ? 32'h13 : _GEN_429; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_431 = 10'h1af == _IFIDIR_T[9:0] ? 32'h13 : _GEN_430; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_432 = 10'h1b0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_431; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_433 = 10'h1b1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_432; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_434 = 10'h1b2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_433; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_435 = 10'h1b3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_434; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_436 = 10'h1b4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_435; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_437 = 10'h1b5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_436; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_438 = 10'h1b6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_437; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_439 = 10'h1b7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_438; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_440 = 10'h1b8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_439; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_441 = 10'h1b9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_440; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_442 = 10'h1ba == _IFIDIR_T[9:0] ? 32'h13 : _GEN_441; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_443 = 10'h1bb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_442; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_444 = 10'h1bc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_443; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_445 = 10'h1bd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_444; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_446 = 10'h1be == _IFIDIR_T[9:0] ? 32'h13 : _GEN_445; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_447 = 10'h1bf == _IFIDIR_T[9:0] ? 32'h13 : _GEN_446; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_448 = 10'h1c0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_447; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_449 = 10'h1c1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_448; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_450 = 10'h1c2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_449; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_451 = 10'h1c3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_450; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_452 = 10'h1c4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_451; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_453 = 10'h1c5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_452; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_454 = 10'h1c6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_453; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_455 = 10'h1c7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_454; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_456 = 10'h1c8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_455; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_457 = 10'h1c9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_456; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_458 = 10'h1ca == _IFIDIR_T[9:0] ? 32'h13 : _GEN_457; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_459 = 10'h1cb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_458; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_460 = 10'h1cc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_459; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_461 = 10'h1cd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_460; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_462 = 10'h1ce == _IFIDIR_T[9:0] ? 32'h13 : _GEN_461; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_463 = 10'h1cf == _IFIDIR_T[9:0] ? 32'h13 : _GEN_462; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_464 = 10'h1d0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_463; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_465 = 10'h1d1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_464; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_466 = 10'h1d2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_465; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_467 = 10'h1d3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_466; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_468 = 10'h1d4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_467; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_469 = 10'h1d5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_468; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_470 = 10'h1d6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_469; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_471 = 10'h1d7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_470; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_472 = 10'h1d8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_471; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_473 = 10'h1d9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_472; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_474 = 10'h1da == _IFIDIR_T[9:0] ? 32'h13 : _GEN_473; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_475 = 10'h1db == _IFIDIR_T[9:0] ? 32'h13 : _GEN_474; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_476 = 10'h1dc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_475; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_477 = 10'h1dd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_476; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_478 = 10'h1de == _IFIDIR_T[9:0] ? 32'h13 : _GEN_477; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_479 = 10'h1df == _IFIDIR_T[9:0] ? 32'h13 : _GEN_478; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_480 = 10'h1e0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_479; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_481 = 10'h1e1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_480; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_482 = 10'h1e2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_481; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_483 = 10'h1e3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_482; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_484 = 10'h1e4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_483; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_485 = 10'h1e5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_484; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_486 = 10'h1e6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_485; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_487 = 10'h1e7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_486; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_488 = 10'h1e8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_487; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_489 = 10'h1e9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_488; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_490 = 10'h1ea == _IFIDIR_T[9:0] ? 32'h13 : _GEN_489; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_491 = 10'h1eb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_490; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_492 = 10'h1ec == _IFIDIR_T[9:0] ? 32'h13 : _GEN_491; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_493 = 10'h1ed == _IFIDIR_T[9:0] ? 32'h13 : _GEN_492; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_494 = 10'h1ee == _IFIDIR_T[9:0] ? 32'h13 : _GEN_493; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_495 = 10'h1ef == _IFIDIR_T[9:0] ? 32'h13 : _GEN_494; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_496 = 10'h1f0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_495; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_497 = 10'h1f1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_496; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_498 = 10'h1f2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_497; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_499 = 10'h1f3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_498; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_500 = 10'h1f4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_499; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_501 = 10'h1f5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_500; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_502 = 10'h1f6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_501; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_503 = 10'h1f7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_502; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_504 = 10'h1f8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_503; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_505 = 10'h1f9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_504; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_506 = 10'h1fa == _IFIDIR_T[9:0] ? 32'h13 : _GEN_505; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_507 = 10'h1fb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_506; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_508 = 10'h1fc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_507; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_509 = 10'h1fd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_508; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_510 = 10'h1fe == _IFIDIR_T[9:0] ? 32'h13 : _GEN_509; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_511 = 10'h1ff == _IFIDIR_T[9:0] ? 32'h13 : _GEN_510; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_512 = 10'h200 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_511; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_513 = 10'h201 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_512; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_514 = 10'h202 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_513; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_515 = 10'h203 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_514; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_516 = 10'h204 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_515; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_517 = 10'h205 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_516; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_518 = 10'h206 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_517; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_519 = 10'h207 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_518; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_520 = 10'h208 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_519; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_521 = 10'h209 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_520; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_522 = 10'h20a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_521; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_523 = 10'h20b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_522; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_524 = 10'h20c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_523; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_525 = 10'h20d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_524; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_526 = 10'h20e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_525; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_527 = 10'h20f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_526; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_528 = 10'h210 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_527; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_529 = 10'h211 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_528; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_530 = 10'h212 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_529; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_531 = 10'h213 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_530; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_532 = 10'h214 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_531; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_533 = 10'h215 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_532; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_534 = 10'h216 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_533; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_535 = 10'h217 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_534; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_536 = 10'h218 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_535; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_537 = 10'h219 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_536; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_538 = 10'h21a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_537; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_539 = 10'h21b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_538; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_540 = 10'h21c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_539; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_541 = 10'h21d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_540; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_542 = 10'h21e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_541; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_543 = 10'h21f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_542; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_544 = 10'h220 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_543; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_545 = 10'h221 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_544; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_546 = 10'h222 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_545; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_547 = 10'h223 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_546; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_548 = 10'h224 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_547; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_549 = 10'h225 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_548; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_550 = 10'h226 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_549; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_551 = 10'h227 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_550; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_552 = 10'h228 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_551; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_553 = 10'h229 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_552; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_554 = 10'h22a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_553; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_555 = 10'h22b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_554; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_556 = 10'h22c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_555; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_557 = 10'h22d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_556; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_558 = 10'h22e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_557; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_559 = 10'h22f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_558; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_560 = 10'h230 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_559; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_561 = 10'h231 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_560; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_562 = 10'h232 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_561; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_563 = 10'h233 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_562; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_564 = 10'h234 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_563; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_565 = 10'h235 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_564; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_566 = 10'h236 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_565; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_567 = 10'h237 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_566; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_568 = 10'h238 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_567; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_569 = 10'h239 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_568; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_570 = 10'h23a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_569; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_571 = 10'h23b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_570; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_572 = 10'h23c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_571; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_573 = 10'h23d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_572; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_574 = 10'h23e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_573; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_575 = 10'h23f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_574; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_576 = 10'h240 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_575; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_577 = 10'h241 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_576; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_578 = 10'h242 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_577; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_579 = 10'h243 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_578; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_580 = 10'h244 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_579; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_581 = 10'h245 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_580; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_582 = 10'h246 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_581; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_583 = 10'h247 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_582; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_584 = 10'h248 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_583; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_585 = 10'h249 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_584; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_586 = 10'h24a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_585; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_587 = 10'h24b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_586; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_588 = 10'h24c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_587; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_589 = 10'h24d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_588; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_590 = 10'h24e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_589; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_591 = 10'h24f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_590; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_592 = 10'h250 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_591; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_593 = 10'h251 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_592; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_594 = 10'h252 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_593; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_595 = 10'h253 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_594; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_596 = 10'h254 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_595; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_597 = 10'h255 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_596; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_598 = 10'h256 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_597; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_599 = 10'h257 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_598; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_600 = 10'h258 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_599; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_601 = 10'h259 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_600; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_602 = 10'h25a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_601; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_603 = 10'h25b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_602; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_604 = 10'h25c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_603; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_605 = 10'h25d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_604; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_606 = 10'h25e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_605; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_607 = 10'h25f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_606; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_608 = 10'h260 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_607; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_609 = 10'h261 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_608; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_610 = 10'h262 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_609; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_611 = 10'h263 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_610; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_612 = 10'h264 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_611; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_613 = 10'h265 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_612; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_614 = 10'h266 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_613; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_615 = 10'h267 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_614; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_616 = 10'h268 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_615; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_617 = 10'h269 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_616; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_618 = 10'h26a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_617; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_619 = 10'h26b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_618; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_620 = 10'h26c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_619; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_621 = 10'h26d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_620; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_622 = 10'h26e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_621; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_623 = 10'h26f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_622; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_624 = 10'h270 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_623; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_625 = 10'h271 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_624; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_626 = 10'h272 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_625; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_627 = 10'h273 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_626; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_628 = 10'h274 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_627; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_629 = 10'h275 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_628; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_630 = 10'h276 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_629; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_631 = 10'h277 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_630; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_632 = 10'h278 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_631; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_633 = 10'h279 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_632; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_634 = 10'h27a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_633; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_635 = 10'h27b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_634; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_636 = 10'h27c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_635; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_637 = 10'h27d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_636; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_638 = 10'h27e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_637; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_639 = 10'h27f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_638; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_640 = 10'h280 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_639; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_641 = 10'h281 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_640; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_642 = 10'h282 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_641; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_643 = 10'h283 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_642; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_644 = 10'h284 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_643; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_645 = 10'h285 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_644; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_646 = 10'h286 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_645; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_647 = 10'h287 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_646; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_648 = 10'h288 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_647; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_649 = 10'h289 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_648; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_650 = 10'h28a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_649; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_651 = 10'h28b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_650; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_652 = 10'h28c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_651; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_653 = 10'h28d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_652; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_654 = 10'h28e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_653; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_655 = 10'h28f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_654; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_656 = 10'h290 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_655; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_657 = 10'h291 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_656; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_658 = 10'h292 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_657; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_659 = 10'h293 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_658; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_660 = 10'h294 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_659; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_661 = 10'h295 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_660; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_662 = 10'h296 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_661; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_663 = 10'h297 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_662; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_664 = 10'h298 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_663; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_665 = 10'h299 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_664; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_666 = 10'h29a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_665; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_667 = 10'h29b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_666; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_668 = 10'h29c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_667; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_669 = 10'h29d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_668; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_670 = 10'h29e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_669; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_671 = 10'h29f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_670; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_672 = 10'h2a0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_671; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_673 = 10'h2a1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_672; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_674 = 10'h2a2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_673; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_675 = 10'h2a3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_674; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_676 = 10'h2a4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_675; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_677 = 10'h2a5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_676; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_678 = 10'h2a6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_677; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_679 = 10'h2a7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_678; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_680 = 10'h2a8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_679; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_681 = 10'h2a9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_680; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_682 = 10'h2aa == _IFIDIR_T[9:0] ? 32'h13 : _GEN_681; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_683 = 10'h2ab == _IFIDIR_T[9:0] ? 32'h13 : _GEN_682; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_684 = 10'h2ac == _IFIDIR_T[9:0] ? 32'h13 : _GEN_683; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_685 = 10'h2ad == _IFIDIR_T[9:0] ? 32'h13 : _GEN_684; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_686 = 10'h2ae == _IFIDIR_T[9:0] ? 32'h13 : _GEN_685; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_687 = 10'h2af == _IFIDIR_T[9:0] ? 32'h13 : _GEN_686; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_688 = 10'h2b0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_687; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_689 = 10'h2b1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_688; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_690 = 10'h2b2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_689; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_691 = 10'h2b3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_690; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_692 = 10'h2b4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_691; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_693 = 10'h2b5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_692; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_694 = 10'h2b6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_693; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_695 = 10'h2b7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_694; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_696 = 10'h2b8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_695; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_697 = 10'h2b9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_696; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_698 = 10'h2ba == _IFIDIR_T[9:0] ? 32'h13 : _GEN_697; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_699 = 10'h2bb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_698; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_700 = 10'h2bc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_699; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_701 = 10'h2bd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_700; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_702 = 10'h2be == _IFIDIR_T[9:0] ? 32'h13 : _GEN_701; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_703 = 10'h2bf == _IFIDIR_T[9:0] ? 32'h13 : _GEN_702; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_704 = 10'h2c0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_703; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_705 = 10'h2c1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_704; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_706 = 10'h2c2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_705; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_707 = 10'h2c3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_706; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_708 = 10'h2c4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_707; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_709 = 10'h2c5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_708; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_710 = 10'h2c6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_709; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_711 = 10'h2c7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_710; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_712 = 10'h2c8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_711; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_713 = 10'h2c9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_712; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_714 = 10'h2ca == _IFIDIR_T[9:0] ? 32'h13 : _GEN_713; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_715 = 10'h2cb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_714; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_716 = 10'h2cc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_715; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_717 = 10'h2cd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_716; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_718 = 10'h2ce == _IFIDIR_T[9:0] ? 32'h13 : _GEN_717; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_719 = 10'h2cf == _IFIDIR_T[9:0] ? 32'h13 : _GEN_718; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_720 = 10'h2d0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_719; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_721 = 10'h2d1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_720; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_722 = 10'h2d2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_721; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_723 = 10'h2d3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_722; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_724 = 10'h2d4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_723; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_725 = 10'h2d5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_724; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_726 = 10'h2d6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_725; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_727 = 10'h2d7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_726; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_728 = 10'h2d8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_727; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_729 = 10'h2d9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_728; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_730 = 10'h2da == _IFIDIR_T[9:0] ? 32'h13 : _GEN_729; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_731 = 10'h2db == _IFIDIR_T[9:0] ? 32'h13 : _GEN_730; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_732 = 10'h2dc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_731; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_733 = 10'h2dd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_732; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_734 = 10'h2de == _IFIDIR_T[9:0] ? 32'h13 : _GEN_733; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_735 = 10'h2df == _IFIDIR_T[9:0] ? 32'h13 : _GEN_734; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_736 = 10'h2e0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_735; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_737 = 10'h2e1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_736; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_738 = 10'h2e2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_737; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_739 = 10'h2e3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_738; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_740 = 10'h2e4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_739; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_741 = 10'h2e5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_740; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_742 = 10'h2e6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_741; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_743 = 10'h2e7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_742; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_744 = 10'h2e8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_743; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_745 = 10'h2e9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_744; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_746 = 10'h2ea == _IFIDIR_T[9:0] ? 32'h13 : _GEN_745; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_747 = 10'h2eb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_746; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_748 = 10'h2ec == _IFIDIR_T[9:0] ? 32'h13 : _GEN_747; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_749 = 10'h2ed == _IFIDIR_T[9:0] ? 32'h13 : _GEN_748; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_750 = 10'h2ee == _IFIDIR_T[9:0] ? 32'h13 : _GEN_749; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_751 = 10'h2ef == _IFIDIR_T[9:0] ? 32'h13 : _GEN_750; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_752 = 10'h2f0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_751; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_753 = 10'h2f1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_752; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_754 = 10'h2f2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_753; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_755 = 10'h2f3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_754; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_756 = 10'h2f4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_755; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_757 = 10'h2f5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_756; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_758 = 10'h2f6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_757; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_759 = 10'h2f7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_758; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_760 = 10'h2f8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_759; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_761 = 10'h2f9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_760; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_762 = 10'h2fa == _IFIDIR_T[9:0] ? 32'h13 : _GEN_761; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_763 = 10'h2fb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_762; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_764 = 10'h2fc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_763; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_765 = 10'h2fd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_764; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_766 = 10'h2fe == _IFIDIR_T[9:0] ? 32'h13 : _GEN_765; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_767 = 10'h2ff == _IFIDIR_T[9:0] ? 32'h13 : _GEN_766; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_768 = 10'h300 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_767; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_769 = 10'h301 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_768; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_770 = 10'h302 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_769; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_771 = 10'h303 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_770; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_772 = 10'h304 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_771; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_773 = 10'h305 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_772; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_774 = 10'h306 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_773; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_775 = 10'h307 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_774; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_776 = 10'h308 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_775; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_777 = 10'h309 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_776; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_778 = 10'h30a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_777; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_779 = 10'h30b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_778; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_780 = 10'h30c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_779; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_781 = 10'h30d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_780; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_782 = 10'h30e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_781; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_783 = 10'h30f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_782; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_784 = 10'h310 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_783; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_785 = 10'h311 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_784; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_786 = 10'h312 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_785; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_787 = 10'h313 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_786; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_788 = 10'h314 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_787; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_789 = 10'h315 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_788; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_790 = 10'h316 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_789; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_791 = 10'h317 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_790; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_792 = 10'h318 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_791; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_793 = 10'h319 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_792; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_794 = 10'h31a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_793; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_795 = 10'h31b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_794; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_796 = 10'h31c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_795; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_797 = 10'h31d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_796; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_798 = 10'h31e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_797; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_799 = 10'h31f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_798; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_800 = 10'h320 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_799; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_801 = 10'h321 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_800; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_802 = 10'h322 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_801; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_803 = 10'h323 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_802; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_804 = 10'h324 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_803; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_805 = 10'h325 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_804; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_806 = 10'h326 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_805; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_807 = 10'h327 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_806; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_808 = 10'h328 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_807; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_809 = 10'h329 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_808; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_810 = 10'h32a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_809; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_811 = 10'h32b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_810; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_812 = 10'h32c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_811; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_813 = 10'h32d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_812; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_814 = 10'h32e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_813; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_815 = 10'h32f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_814; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_816 = 10'h330 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_815; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_817 = 10'h331 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_816; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_818 = 10'h332 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_817; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_819 = 10'h333 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_818; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_820 = 10'h334 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_819; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_821 = 10'h335 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_820; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_822 = 10'h336 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_821; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_823 = 10'h337 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_822; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_824 = 10'h338 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_823; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_825 = 10'h339 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_824; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_826 = 10'h33a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_825; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_827 = 10'h33b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_826; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_828 = 10'h33c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_827; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_829 = 10'h33d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_828; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_830 = 10'h33e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_829; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_831 = 10'h33f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_830; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_832 = 10'h340 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_831; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_833 = 10'h341 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_832; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_834 = 10'h342 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_833; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_835 = 10'h343 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_834; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_836 = 10'h344 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_835; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_837 = 10'h345 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_836; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_838 = 10'h346 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_837; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_839 = 10'h347 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_838; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_840 = 10'h348 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_839; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_841 = 10'h349 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_840; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_842 = 10'h34a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_841; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_843 = 10'h34b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_842; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_844 = 10'h34c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_843; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_845 = 10'h34d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_844; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_846 = 10'h34e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_845; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_847 = 10'h34f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_846; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_848 = 10'h350 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_847; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_849 = 10'h351 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_848; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_850 = 10'h352 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_849; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_851 = 10'h353 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_850; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_852 = 10'h354 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_851; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_853 = 10'h355 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_852; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_854 = 10'h356 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_853; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_855 = 10'h357 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_854; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_856 = 10'h358 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_855; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_857 = 10'h359 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_856; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_858 = 10'h35a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_857; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_859 = 10'h35b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_858; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_860 = 10'h35c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_859; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_861 = 10'h35d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_860; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_862 = 10'h35e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_861; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_863 = 10'h35f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_862; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_864 = 10'h360 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_863; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_865 = 10'h361 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_864; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_866 = 10'h362 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_865; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_867 = 10'h363 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_866; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_868 = 10'h364 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_867; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_869 = 10'h365 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_868; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_870 = 10'h366 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_869; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_871 = 10'h367 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_870; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_872 = 10'h368 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_871; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_873 = 10'h369 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_872; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_874 = 10'h36a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_873; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_875 = 10'h36b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_874; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_876 = 10'h36c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_875; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_877 = 10'h36d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_876; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_878 = 10'h36e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_877; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_879 = 10'h36f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_878; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_880 = 10'h370 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_879; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_881 = 10'h371 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_880; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_882 = 10'h372 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_881; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_883 = 10'h373 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_882; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_884 = 10'h374 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_883; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_885 = 10'h375 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_884; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_886 = 10'h376 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_885; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_887 = 10'h377 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_886; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_888 = 10'h378 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_887; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_889 = 10'h379 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_888; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_890 = 10'h37a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_889; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_891 = 10'h37b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_890; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_892 = 10'h37c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_891; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_893 = 10'h37d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_892; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_894 = 10'h37e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_893; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_895 = 10'h37f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_894; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_896 = 10'h380 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_895; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_897 = 10'h381 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_896; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_898 = 10'h382 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_897; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_899 = 10'h383 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_898; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_900 = 10'h384 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_899; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_901 = 10'h385 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_900; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_902 = 10'h386 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_901; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_903 = 10'h387 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_902; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_904 = 10'h388 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_903; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_905 = 10'h389 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_904; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_906 = 10'h38a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_905; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_907 = 10'h38b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_906; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_908 = 10'h38c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_907; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_909 = 10'h38d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_908; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_910 = 10'h38e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_909; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_911 = 10'h38f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_910; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_912 = 10'h390 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_911; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_913 = 10'h391 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_912; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_914 = 10'h392 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_913; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_915 = 10'h393 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_914; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_916 = 10'h394 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_915; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_917 = 10'h395 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_916; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_918 = 10'h396 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_917; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_919 = 10'h397 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_918; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_920 = 10'h398 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_919; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_921 = 10'h399 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_920; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_922 = 10'h39a == _IFIDIR_T[9:0] ? 32'h13 : _GEN_921; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_923 = 10'h39b == _IFIDIR_T[9:0] ? 32'h13 : _GEN_922; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_924 = 10'h39c == _IFIDIR_T[9:0] ? 32'h13 : _GEN_923; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_925 = 10'h39d == _IFIDIR_T[9:0] ? 32'h13 : _GEN_924; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_926 = 10'h39e == _IFIDIR_T[9:0] ? 32'h13 : _GEN_925; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_927 = 10'h39f == _IFIDIR_T[9:0] ? 32'h13 : _GEN_926; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_928 = 10'h3a0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_927; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_929 = 10'h3a1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_928; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_930 = 10'h3a2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_929; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_931 = 10'h3a3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_930; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_932 = 10'h3a4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_931; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_933 = 10'h3a5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_932; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_934 = 10'h3a6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_933; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_935 = 10'h3a7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_934; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_936 = 10'h3a8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_935; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_937 = 10'h3a9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_936; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_938 = 10'h3aa == _IFIDIR_T[9:0] ? 32'h13 : _GEN_937; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_939 = 10'h3ab == _IFIDIR_T[9:0] ? 32'h13 : _GEN_938; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_940 = 10'h3ac == _IFIDIR_T[9:0] ? 32'h13 : _GEN_939; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_941 = 10'h3ad == _IFIDIR_T[9:0] ? 32'h13 : _GEN_940; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_942 = 10'h3ae == _IFIDIR_T[9:0] ? 32'h13 : _GEN_941; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_943 = 10'h3af == _IFIDIR_T[9:0] ? 32'h13 : _GEN_942; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_944 = 10'h3b0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_943; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_945 = 10'h3b1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_944; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_946 = 10'h3b2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_945; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_947 = 10'h3b3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_946; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_948 = 10'h3b4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_947; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_949 = 10'h3b5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_948; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_950 = 10'h3b6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_949; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_951 = 10'h3b7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_950; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_952 = 10'h3b8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_951; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_953 = 10'h3b9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_952; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_954 = 10'h3ba == _IFIDIR_T[9:0] ? 32'h13 : _GEN_953; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_955 = 10'h3bb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_954; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_956 = 10'h3bc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_955; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_957 = 10'h3bd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_956; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_958 = 10'h3be == _IFIDIR_T[9:0] ? 32'h13 : _GEN_957; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_959 = 10'h3bf == _IFIDIR_T[9:0] ? 32'h13 : _GEN_958; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_960 = 10'h3c0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_959; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_961 = 10'h3c1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_960; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_962 = 10'h3c2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_961; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_963 = 10'h3c3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_962; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_964 = 10'h3c4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_963; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_965 = 10'h3c5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_964; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_966 = 10'h3c6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_965; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_967 = 10'h3c7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_966; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_968 = 10'h3c8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_967; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_969 = 10'h3c9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_968; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_970 = 10'h3ca == _IFIDIR_T[9:0] ? 32'h13 : _GEN_969; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_971 = 10'h3cb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_970; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_972 = 10'h3cc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_971; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_973 = 10'h3cd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_972; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_974 = 10'h3ce == _IFIDIR_T[9:0] ? 32'h13 : _GEN_973; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_975 = 10'h3cf == _IFIDIR_T[9:0] ? 32'h13 : _GEN_974; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_976 = 10'h3d0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_975; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_977 = 10'h3d1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_976; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_978 = 10'h3d2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_977; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_979 = 10'h3d3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_978; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_980 = 10'h3d4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_979; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_981 = 10'h3d5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_980; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_982 = 10'h3d6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_981; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_983 = 10'h3d7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_982; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_984 = 10'h3d8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_983; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_985 = 10'h3d9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_984; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_986 = 10'h3da == _IFIDIR_T[9:0] ? 32'h13 : _GEN_985; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_987 = 10'h3db == _IFIDIR_T[9:0] ? 32'h13 : _GEN_986; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_988 = 10'h3dc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_987; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_989 = 10'h3dd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_988; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_990 = 10'h3de == _IFIDIR_T[9:0] ? 32'h13 : _GEN_989; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_991 = 10'h3df == _IFIDIR_T[9:0] ? 32'h13 : _GEN_990; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_992 = 10'h3e0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_991; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_993 = 10'h3e1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_992; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_994 = 10'h3e2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_993; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_995 = 10'h3e3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_994; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_996 = 10'h3e4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_995; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_997 = 10'h3e5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_996; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_998 = 10'h3e6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_997; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_999 = 10'h3e7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_998; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1000 = 10'h3e8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_999; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1001 = 10'h3e9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1000; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1002 = 10'h3ea == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1001; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1003 = 10'h3eb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1002; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1004 = 10'h3ec == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1003; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1005 = 10'h3ed == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1004; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1006 = 10'h3ee == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1005; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1007 = 10'h3ef == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1006; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1008 = 10'h3f0 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1007; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1009 = 10'h3f1 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1008; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1010 = 10'h3f2 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1009; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1011 = 10'h3f3 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1010; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1012 = 10'h3f4 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1011; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1013 = 10'h3f5 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1012; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1014 = 10'h3f6 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1013; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1015 = 10'h3f7 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1014; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1016 = 10'h3f8 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1015; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1017 = 10'h3f9 == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1016; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1018 = 10'h3fa == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1017; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1019 = 10'h3fb == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1018; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1020 = 10'h3fc == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1019; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1021 = 10'h3fd == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1020; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1022 = 10'h3fe == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1021; // @[cpu.scala 141:{16,16}]
  wire [31:0] _GEN_1023 = 10'h3ff == _IFIDIR_T[9:0] ? 32'h13 : _GEN_1022; // @[cpu.scala 141:{16,16}]
  wire [63:0] _PC_T_1 = PC + 64'h4; // @[cpu.scala 142:18]
  wire [12:0] _branchTarget_T_5 = {IFIDIR[31],1'h0,IFIDIR[30:25],IFIDIR[11:7]}; // @[cpu.scala 151:11]
  wire [63:0] _GEN_7388 = {{51{_branchTarget_T_5[12]}},_branchTarget_T_5}; // @[cpu.scala 146:42]
  wire [63:0] branchTarget = $signed(CurPC) + $signed(_GEN_7388); // @[cpu.scala 151:19]
  wire [11:0] _EXMEMALUOut_T_2 = IDEXIR[31:20]; // @[cpu.scala 199:53]
  wire [63:0] _GEN_7389 = {{52{_EXMEMALUOut_T_2[11]}},_EXMEMALUOut_T_2}; // @[cpu.scala 199:36]
  wire [63:0] _EXMEMALUOut_T_6 = $signed(IDEXA) + $signed(_GEN_7389); // @[cpu.scala 199:61]
  wire [11:0] _EXMEMALUOut_T_11 = {IDEXIR[31:25],IDEXrd}; // @[cpu.scala 204:9]
  wire [63:0] _GEN_7390 = {{52{_EXMEMALUOut_T_11[11]}},_EXMEMALUOut_T_11}; // @[cpu.scala 201:36]
  wire [63:0] _EXMEMALUOut_T_15 = $signed(IDEXA) + $signed(_GEN_7390); // @[cpu.scala 204:17]
  wire [31:0] _GEN_1118 = 10'h1 == EXMEMALUOut[9:0] ? DMemory_1 : DMemory_0; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1119 = 10'h2 == EXMEMALUOut[9:0] ? DMemory_2 : _GEN_1118; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1120 = 10'h3 == EXMEMALUOut[9:0] ? DMemory_3 : _GEN_1119; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1121 = 10'h4 == EXMEMALUOut[9:0] ? DMemory_4 : _GEN_1120; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1122 = 10'h5 == EXMEMALUOut[9:0] ? DMemory_5 : _GEN_1121; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1123 = 10'h6 == EXMEMALUOut[9:0] ? DMemory_6 : _GEN_1122; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1124 = 10'h7 == EXMEMALUOut[9:0] ? DMemory_7 : _GEN_1123; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1125 = 10'h8 == EXMEMALUOut[9:0] ? DMemory_8 : _GEN_1124; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1126 = 10'h9 == EXMEMALUOut[9:0] ? DMemory_9 : _GEN_1125; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1127 = 10'ha == EXMEMALUOut[9:0] ? DMemory_10 : _GEN_1126; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1128 = 10'hb == EXMEMALUOut[9:0] ? DMemory_11 : _GEN_1127; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1129 = 10'hc == EXMEMALUOut[9:0] ? DMemory_12 : _GEN_1128; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1130 = 10'hd == EXMEMALUOut[9:0] ? DMemory_13 : _GEN_1129; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1131 = 10'he == EXMEMALUOut[9:0] ? DMemory_14 : _GEN_1130; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1132 = 10'hf == EXMEMALUOut[9:0] ? DMemory_15 : _GEN_1131; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1133 = 10'h10 == EXMEMALUOut[9:0] ? DMemory_16 : _GEN_1132; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1134 = 10'h11 == EXMEMALUOut[9:0] ? DMemory_17 : _GEN_1133; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1135 = 10'h12 == EXMEMALUOut[9:0] ? DMemory_18 : _GEN_1134; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1136 = 10'h13 == EXMEMALUOut[9:0] ? DMemory_19 : _GEN_1135; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1137 = 10'h14 == EXMEMALUOut[9:0] ? DMemory_20 : _GEN_1136; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1138 = 10'h15 == EXMEMALUOut[9:0] ? DMemory_21 : _GEN_1137; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1139 = 10'h16 == EXMEMALUOut[9:0] ? DMemory_22 : _GEN_1138; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1140 = 10'h17 == EXMEMALUOut[9:0] ? DMemory_23 : _GEN_1139; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1141 = 10'h18 == EXMEMALUOut[9:0] ? DMemory_24 : _GEN_1140; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1142 = 10'h19 == EXMEMALUOut[9:0] ? DMemory_25 : _GEN_1141; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1143 = 10'h1a == EXMEMALUOut[9:0] ? DMemory_26 : _GEN_1142; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1144 = 10'h1b == EXMEMALUOut[9:0] ? DMemory_27 : _GEN_1143; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1145 = 10'h1c == EXMEMALUOut[9:0] ? DMemory_28 : _GEN_1144; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1146 = 10'h1d == EXMEMALUOut[9:0] ? DMemory_29 : _GEN_1145; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1147 = 10'h1e == EXMEMALUOut[9:0] ? DMemory_30 : _GEN_1146; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1148 = 10'h1f == EXMEMALUOut[9:0] ? DMemory_31 : _GEN_1147; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1149 = 10'h20 == EXMEMALUOut[9:0] ? DMemory_32 : _GEN_1148; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1150 = 10'h21 == EXMEMALUOut[9:0] ? DMemory_33 : _GEN_1149; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1151 = 10'h22 == EXMEMALUOut[9:0] ? DMemory_34 : _GEN_1150; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1152 = 10'h23 == EXMEMALUOut[9:0] ? DMemory_35 : _GEN_1151; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1153 = 10'h24 == EXMEMALUOut[9:0] ? DMemory_36 : _GEN_1152; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1154 = 10'h25 == EXMEMALUOut[9:0] ? DMemory_37 : _GEN_1153; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1155 = 10'h26 == EXMEMALUOut[9:0] ? DMemory_38 : _GEN_1154; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1156 = 10'h27 == EXMEMALUOut[9:0] ? DMemory_39 : _GEN_1155; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1157 = 10'h28 == EXMEMALUOut[9:0] ? DMemory_40 : _GEN_1156; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1158 = 10'h29 == EXMEMALUOut[9:0] ? DMemory_41 : _GEN_1157; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1159 = 10'h2a == EXMEMALUOut[9:0] ? DMemory_42 : _GEN_1158; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1160 = 10'h2b == EXMEMALUOut[9:0] ? DMemory_43 : _GEN_1159; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1161 = 10'h2c == EXMEMALUOut[9:0] ? DMemory_44 : _GEN_1160; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1162 = 10'h2d == EXMEMALUOut[9:0] ? DMemory_45 : _GEN_1161; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1163 = 10'h2e == EXMEMALUOut[9:0] ? DMemory_46 : _GEN_1162; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1164 = 10'h2f == EXMEMALUOut[9:0] ? DMemory_47 : _GEN_1163; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1165 = 10'h30 == EXMEMALUOut[9:0] ? DMemory_48 : _GEN_1164; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1166 = 10'h31 == EXMEMALUOut[9:0] ? DMemory_49 : _GEN_1165; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1167 = 10'h32 == EXMEMALUOut[9:0] ? DMemory_50 : _GEN_1166; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1168 = 10'h33 == EXMEMALUOut[9:0] ? DMemory_51 : _GEN_1167; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1169 = 10'h34 == EXMEMALUOut[9:0] ? DMemory_52 : _GEN_1168; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1170 = 10'h35 == EXMEMALUOut[9:0] ? DMemory_53 : _GEN_1169; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1171 = 10'h36 == EXMEMALUOut[9:0] ? DMemory_54 : _GEN_1170; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1172 = 10'h37 == EXMEMALUOut[9:0] ? DMemory_55 : _GEN_1171; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1173 = 10'h38 == EXMEMALUOut[9:0] ? DMemory_56 : _GEN_1172; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1174 = 10'h39 == EXMEMALUOut[9:0] ? DMemory_57 : _GEN_1173; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1175 = 10'h3a == EXMEMALUOut[9:0] ? DMemory_58 : _GEN_1174; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1176 = 10'h3b == EXMEMALUOut[9:0] ? DMemory_59 : _GEN_1175; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1177 = 10'h3c == EXMEMALUOut[9:0] ? DMemory_60 : _GEN_1176; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1178 = 10'h3d == EXMEMALUOut[9:0] ? DMemory_61 : _GEN_1177; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1179 = 10'h3e == EXMEMALUOut[9:0] ? DMemory_62 : _GEN_1178; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1180 = 10'h3f == EXMEMALUOut[9:0] ? DMemory_63 : _GEN_1179; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1181 = 10'h40 == EXMEMALUOut[9:0] ? DMemory_64 : _GEN_1180; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1182 = 10'h41 == EXMEMALUOut[9:0] ? DMemory_65 : _GEN_1181; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1183 = 10'h42 == EXMEMALUOut[9:0] ? DMemory_66 : _GEN_1182; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1184 = 10'h43 == EXMEMALUOut[9:0] ? DMemory_67 : _GEN_1183; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1185 = 10'h44 == EXMEMALUOut[9:0] ? DMemory_68 : _GEN_1184; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1186 = 10'h45 == EXMEMALUOut[9:0] ? DMemory_69 : _GEN_1185; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1187 = 10'h46 == EXMEMALUOut[9:0] ? DMemory_70 : _GEN_1186; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1188 = 10'h47 == EXMEMALUOut[9:0] ? DMemory_71 : _GEN_1187; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1189 = 10'h48 == EXMEMALUOut[9:0] ? DMemory_72 : _GEN_1188; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1190 = 10'h49 == EXMEMALUOut[9:0] ? DMemory_73 : _GEN_1189; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1191 = 10'h4a == EXMEMALUOut[9:0] ? DMemory_74 : _GEN_1190; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1192 = 10'h4b == EXMEMALUOut[9:0] ? DMemory_75 : _GEN_1191; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1193 = 10'h4c == EXMEMALUOut[9:0] ? DMemory_76 : _GEN_1192; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1194 = 10'h4d == EXMEMALUOut[9:0] ? DMemory_77 : _GEN_1193; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1195 = 10'h4e == EXMEMALUOut[9:0] ? DMemory_78 : _GEN_1194; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1196 = 10'h4f == EXMEMALUOut[9:0] ? DMemory_79 : _GEN_1195; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1197 = 10'h50 == EXMEMALUOut[9:0] ? DMemory_80 : _GEN_1196; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1198 = 10'h51 == EXMEMALUOut[9:0] ? DMemory_81 : _GEN_1197; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1199 = 10'h52 == EXMEMALUOut[9:0] ? DMemory_82 : _GEN_1198; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1200 = 10'h53 == EXMEMALUOut[9:0] ? DMemory_83 : _GEN_1199; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1201 = 10'h54 == EXMEMALUOut[9:0] ? DMemory_84 : _GEN_1200; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1202 = 10'h55 == EXMEMALUOut[9:0] ? DMemory_85 : _GEN_1201; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1203 = 10'h56 == EXMEMALUOut[9:0] ? DMemory_86 : _GEN_1202; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1204 = 10'h57 == EXMEMALUOut[9:0] ? DMemory_87 : _GEN_1203; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1205 = 10'h58 == EXMEMALUOut[9:0] ? DMemory_88 : _GEN_1204; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1206 = 10'h59 == EXMEMALUOut[9:0] ? DMemory_89 : _GEN_1205; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1207 = 10'h5a == EXMEMALUOut[9:0] ? DMemory_90 : _GEN_1206; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1208 = 10'h5b == EXMEMALUOut[9:0] ? DMemory_91 : _GEN_1207; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1209 = 10'h5c == EXMEMALUOut[9:0] ? DMemory_92 : _GEN_1208; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1210 = 10'h5d == EXMEMALUOut[9:0] ? DMemory_93 : _GEN_1209; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1211 = 10'h5e == EXMEMALUOut[9:0] ? DMemory_94 : _GEN_1210; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1212 = 10'h5f == EXMEMALUOut[9:0] ? DMemory_95 : _GEN_1211; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1213 = 10'h60 == EXMEMALUOut[9:0] ? DMemory_96 : _GEN_1212; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1214 = 10'h61 == EXMEMALUOut[9:0] ? DMemory_97 : _GEN_1213; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1215 = 10'h62 == EXMEMALUOut[9:0] ? DMemory_98 : _GEN_1214; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1216 = 10'h63 == EXMEMALUOut[9:0] ? DMemory_99 : _GEN_1215; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1217 = 10'h64 == EXMEMALUOut[9:0] ? DMemory_100 : _GEN_1216; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1218 = 10'h65 == EXMEMALUOut[9:0] ? DMemory_101 : _GEN_1217; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1219 = 10'h66 == EXMEMALUOut[9:0] ? DMemory_102 : _GEN_1218; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1220 = 10'h67 == EXMEMALUOut[9:0] ? DMemory_103 : _GEN_1219; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1221 = 10'h68 == EXMEMALUOut[9:0] ? DMemory_104 : _GEN_1220; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1222 = 10'h69 == EXMEMALUOut[9:0] ? DMemory_105 : _GEN_1221; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1223 = 10'h6a == EXMEMALUOut[9:0] ? DMemory_106 : _GEN_1222; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1224 = 10'h6b == EXMEMALUOut[9:0] ? DMemory_107 : _GEN_1223; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1225 = 10'h6c == EXMEMALUOut[9:0] ? DMemory_108 : _GEN_1224; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1226 = 10'h6d == EXMEMALUOut[9:0] ? DMemory_109 : _GEN_1225; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1227 = 10'h6e == EXMEMALUOut[9:0] ? DMemory_110 : _GEN_1226; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1228 = 10'h6f == EXMEMALUOut[9:0] ? DMemory_111 : _GEN_1227; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1229 = 10'h70 == EXMEMALUOut[9:0] ? DMemory_112 : _GEN_1228; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1230 = 10'h71 == EXMEMALUOut[9:0] ? DMemory_113 : _GEN_1229; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1231 = 10'h72 == EXMEMALUOut[9:0] ? DMemory_114 : _GEN_1230; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1232 = 10'h73 == EXMEMALUOut[9:0] ? DMemory_115 : _GEN_1231; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1233 = 10'h74 == EXMEMALUOut[9:0] ? DMemory_116 : _GEN_1232; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1234 = 10'h75 == EXMEMALUOut[9:0] ? DMemory_117 : _GEN_1233; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1235 = 10'h76 == EXMEMALUOut[9:0] ? DMemory_118 : _GEN_1234; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1236 = 10'h77 == EXMEMALUOut[9:0] ? DMemory_119 : _GEN_1235; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1237 = 10'h78 == EXMEMALUOut[9:0] ? DMemory_120 : _GEN_1236; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1238 = 10'h79 == EXMEMALUOut[9:0] ? DMemory_121 : _GEN_1237; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1239 = 10'h7a == EXMEMALUOut[9:0] ? DMemory_122 : _GEN_1238; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1240 = 10'h7b == EXMEMALUOut[9:0] ? DMemory_123 : _GEN_1239; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1241 = 10'h7c == EXMEMALUOut[9:0] ? DMemory_124 : _GEN_1240; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1242 = 10'h7d == EXMEMALUOut[9:0] ? DMemory_125 : _GEN_1241; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1243 = 10'h7e == EXMEMALUOut[9:0] ? DMemory_126 : _GEN_1242; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1244 = 10'h7f == EXMEMALUOut[9:0] ? DMemory_127 : _GEN_1243; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1245 = 10'h80 == EXMEMALUOut[9:0] ? DMemory_128 : _GEN_1244; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1246 = 10'h81 == EXMEMALUOut[9:0] ? DMemory_129 : _GEN_1245; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1247 = 10'h82 == EXMEMALUOut[9:0] ? DMemory_130 : _GEN_1246; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1248 = 10'h83 == EXMEMALUOut[9:0] ? DMemory_131 : _GEN_1247; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1249 = 10'h84 == EXMEMALUOut[9:0] ? DMemory_132 : _GEN_1248; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1250 = 10'h85 == EXMEMALUOut[9:0] ? DMemory_133 : _GEN_1249; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1251 = 10'h86 == EXMEMALUOut[9:0] ? DMemory_134 : _GEN_1250; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1252 = 10'h87 == EXMEMALUOut[9:0] ? DMemory_135 : _GEN_1251; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1253 = 10'h88 == EXMEMALUOut[9:0] ? DMemory_136 : _GEN_1252; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1254 = 10'h89 == EXMEMALUOut[9:0] ? DMemory_137 : _GEN_1253; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1255 = 10'h8a == EXMEMALUOut[9:0] ? DMemory_138 : _GEN_1254; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1256 = 10'h8b == EXMEMALUOut[9:0] ? DMemory_139 : _GEN_1255; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1257 = 10'h8c == EXMEMALUOut[9:0] ? DMemory_140 : _GEN_1256; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1258 = 10'h8d == EXMEMALUOut[9:0] ? DMemory_141 : _GEN_1257; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1259 = 10'h8e == EXMEMALUOut[9:0] ? DMemory_142 : _GEN_1258; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1260 = 10'h8f == EXMEMALUOut[9:0] ? DMemory_143 : _GEN_1259; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1261 = 10'h90 == EXMEMALUOut[9:0] ? DMemory_144 : _GEN_1260; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1262 = 10'h91 == EXMEMALUOut[9:0] ? DMemory_145 : _GEN_1261; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1263 = 10'h92 == EXMEMALUOut[9:0] ? DMemory_146 : _GEN_1262; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1264 = 10'h93 == EXMEMALUOut[9:0] ? DMemory_147 : _GEN_1263; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1265 = 10'h94 == EXMEMALUOut[9:0] ? DMemory_148 : _GEN_1264; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1266 = 10'h95 == EXMEMALUOut[9:0] ? DMemory_149 : _GEN_1265; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1267 = 10'h96 == EXMEMALUOut[9:0] ? DMemory_150 : _GEN_1266; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1268 = 10'h97 == EXMEMALUOut[9:0] ? DMemory_151 : _GEN_1267; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1269 = 10'h98 == EXMEMALUOut[9:0] ? DMemory_152 : _GEN_1268; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1270 = 10'h99 == EXMEMALUOut[9:0] ? DMemory_153 : _GEN_1269; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1271 = 10'h9a == EXMEMALUOut[9:0] ? DMemory_154 : _GEN_1270; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1272 = 10'h9b == EXMEMALUOut[9:0] ? DMemory_155 : _GEN_1271; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1273 = 10'h9c == EXMEMALUOut[9:0] ? DMemory_156 : _GEN_1272; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1274 = 10'h9d == EXMEMALUOut[9:0] ? DMemory_157 : _GEN_1273; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1275 = 10'h9e == EXMEMALUOut[9:0] ? DMemory_158 : _GEN_1274; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1276 = 10'h9f == EXMEMALUOut[9:0] ? DMemory_159 : _GEN_1275; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1277 = 10'ha0 == EXMEMALUOut[9:0] ? DMemory_160 : _GEN_1276; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1278 = 10'ha1 == EXMEMALUOut[9:0] ? DMemory_161 : _GEN_1277; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1279 = 10'ha2 == EXMEMALUOut[9:0] ? DMemory_162 : _GEN_1278; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1280 = 10'ha3 == EXMEMALUOut[9:0] ? DMemory_163 : _GEN_1279; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1281 = 10'ha4 == EXMEMALUOut[9:0] ? DMemory_164 : _GEN_1280; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1282 = 10'ha5 == EXMEMALUOut[9:0] ? DMemory_165 : _GEN_1281; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1283 = 10'ha6 == EXMEMALUOut[9:0] ? DMemory_166 : _GEN_1282; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1284 = 10'ha7 == EXMEMALUOut[9:0] ? DMemory_167 : _GEN_1283; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1285 = 10'ha8 == EXMEMALUOut[9:0] ? DMemory_168 : _GEN_1284; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1286 = 10'ha9 == EXMEMALUOut[9:0] ? DMemory_169 : _GEN_1285; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1287 = 10'haa == EXMEMALUOut[9:0] ? DMemory_170 : _GEN_1286; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1288 = 10'hab == EXMEMALUOut[9:0] ? DMemory_171 : _GEN_1287; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1289 = 10'hac == EXMEMALUOut[9:0] ? DMemory_172 : _GEN_1288; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1290 = 10'had == EXMEMALUOut[9:0] ? DMemory_173 : _GEN_1289; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1291 = 10'hae == EXMEMALUOut[9:0] ? DMemory_174 : _GEN_1290; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1292 = 10'haf == EXMEMALUOut[9:0] ? DMemory_175 : _GEN_1291; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1293 = 10'hb0 == EXMEMALUOut[9:0] ? DMemory_176 : _GEN_1292; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1294 = 10'hb1 == EXMEMALUOut[9:0] ? DMemory_177 : _GEN_1293; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1295 = 10'hb2 == EXMEMALUOut[9:0] ? DMemory_178 : _GEN_1294; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1296 = 10'hb3 == EXMEMALUOut[9:0] ? DMemory_179 : _GEN_1295; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1297 = 10'hb4 == EXMEMALUOut[9:0] ? DMemory_180 : _GEN_1296; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1298 = 10'hb5 == EXMEMALUOut[9:0] ? DMemory_181 : _GEN_1297; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1299 = 10'hb6 == EXMEMALUOut[9:0] ? DMemory_182 : _GEN_1298; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1300 = 10'hb7 == EXMEMALUOut[9:0] ? DMemory_183 : _GEN_1299; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1301 = 10'hb8 == EXMEMALUOut[9:0] ? DMemory_184 : _GEN_1300; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1302 = 10'hb9 == EXMEMALUOut[9:0] ? DMemory_185 : _GEN_1301; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1303 = 10'hba == EXMEMALUOut[9:0] ? DMemory_186 : _GEN_1302; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1304 = 10'hbb == EXMEMALUOut[9:0] ? DMemory_187 : _GEN_1303; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1305 = 10'hbc == EXMEMALUOut[9:0] ? DMemory_188 : _GEN_1304; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1306 = 10'hbd == EXMEMALUOut[9:0] ? DMemory_189 : _GEN_1305; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1307 = 10'hbe == EXMEMALUOut[9:0] ? DMemory_190 : _GEN_1306; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1308 = 10'hbf == EXMEMALUOut[9:0] ? DMemory_191 : _GEN_1307; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1309 = 10'hc0 == EXMEMALUOut[9:0] ? DMemory_192 : _GEN_1308; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1310 = 10'hc1 == EXMEMALUOut[9:0] ? DMemory_193 : _GEN_1309; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1311 = 10'hc2 == EXMEMALUOut[9:0] ? DMemory_194 : _GEN_1310; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1312 = 10'hc3 == EXMEMALUOut[9:0] ? DMemory_195 : _GEN_1311; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1313 = 10'hc4 == EXMEMALUOut[9:0] ? DMemory_196 : _GEN_1312; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1314 = 10'hc5 == EXMEMALUOut[9:0] ? DMemory_197 : _GEN_1313; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1315 = 10'hc6 == EXMEMALUOut[9:0] ? DMemory_198 : _GEN_1314; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1316 = 10'hc7 == EXMEMALUOut[9:0] ? DMemory_199 : _GEN_1315; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1317 = 10'hc8 == EXMEMALUOut[9:0] ? DMemory_200 : _GEN_1316; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1318 = 10'hc9 == EXMEMALUOut[9:0] ? DMemory_201 : _GEN_1317; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1319 = 10'hca == EXMEMALUOut[9:0] ? DMemory_202 : _GEN_1318; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1320 = 10'hcb == EXMEMALUOut[9:0] ? DMemory_203 : _GEN_1319; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1321 = 10'hcc == EXMEMALUOut[9:0] ? DMemory_204 : _GEN_1320; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1322 = 10'hcd == EXMEMALUOut[9:0] ? DMemory_205 : _GEN_1321; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1323 = 10'hce == EXMEMALUOut[9:0] ? DMemory_206 : _GEN_1322; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1324 = 10'hcf == EXMEMALUOut[9:0] ? DMemory_207 : _GEN_1323; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1325 = 10'hd0 == EXMEMALUOut[9:0] ? DMemory_208 : _GEN_1324; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1326 = 10'hd1 == EXMEMALUOut[9:0] ? DMemory_209 : _GEN_1325; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1327 = 10'hd2 == EXMEMALUOut[9:0] ? DMemory_210 : _GEN_1326; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1328 = 10'hd3 == EXMEMALUOut[9:0] ? DMemory_211 : _GEN_1327; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1329 = 10'hd4 == EXMEMALUOut[9:0] ? DMemory_212 : _GEN_1328; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1330 = 10'hd5 == EXMEMALUOut[9:0] ? DMemory_213 : _GEN_1329; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1331 = 10'hd6 == EXMEMALUOut[9:0] ? DMemory_214 : _GEN_1330; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1332 = 10'hd7 == EXMEMALUOut[9:0] ? DMemory_215 : _GEN_1331; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1333 = 10'hd8 == EXMEMALUOut[9:0] ? DMemory_216 : _GEN_1332; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1334 = 10'hd9 == EXMEMALUOut[9:0] ? DMemory_217 : _GEN_1333; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1335 = 10'hda == EXMEMALUOut[9:0] ? DMemory_218 : _GEN_1334; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1336 = 10'hdb == EXMEMALUOut[9:0] ? DMemory_219 : _GEN_1335; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1337 = 10'hdc == EXMEMALUOut[9:0] ? DMemory_220 : _GEN_1336; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1338 = 10'hdd == EXMEMALUOut[9:0] ? DMemory_221 : _GEN_1337; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1339 = 10'hde == EXMEMALUOut[9:0] ? DMemory_222 : _GEN_1338; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1340 = 10'hdf == EXMEMALUOut[9:0] ? DMemory_223 : _GEN_1339; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1341 = 10'he0 == EXMEMALUOut[9:0] ? DMemory_224 : _GEN_1340; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1342 = 10'he1 == EXMEMALUOut[9:0] ? DMemory_225 : _GEN_1341; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1343 = 10'he2 == EXMEMALUOut[9:0] ? DMemory_226 : _GEN_1342; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1344 = 10'he3 == EXMEMALUOut[9:0] ? DMemory_227 : _GEN_1343; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1345 = 10'he4 == EXMEMALUOut[9:0] ? DMemory_228 : _GEN_1344; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1346 = 10'he5 == EXMEMALUOut[9:0] ? DMemory_229 : _GEN_1345; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1347 = 10'he6 == EXMEMALUOut[9:0] ? DMemory_230 : _GEN_1346; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1348 = 10'he7 == EXMEMALUOut[9:0] ? DMemory_231 : _GEN_1347; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1349 = 10'he8 == EXMEMALUOut[9:0] ? DMemory_232 : _GEN_1348; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1350 = 10'he9 == EXMEMALUOut[9:0] ? DMemory_233 : _GEN_1349; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1351 = 10'hea == EXMEMALUOut[9:0] ? DMemory_234 : _GEN_1350; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1352 = 10'heb == EXMEMALUOut[9:0] ? DMemory_235 : _GEN_1351; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1353 = 10'hec == EXMEMALUOut[9:0] ? DMemory_236 : _GEN_1352; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1354 = 10'hed == EXMEMALUOut[9:0] ? DMemory_237 : _GEN_1353; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1355 = 10'hee == EXMEMALUOut[9:0] ? DMemory_238 : _GEN_1354; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1356 = 10'hef == EXMEMALUOut[9:0] ? DMemory_239 : _GEN_1355; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1357 = 10'hf0 == EXMEMALUOut[9:0] ? DMemory_240 : _GEN_1356; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1358 = 10'hf1 == EXMEMALUOut[9:0] ? DMemory_241 : _GEN_1357; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1359 = 10'hf2 == EXMEMALUOut[9:0] ? DMemory_242 : _GEN_1358; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1360 = 10'hf3 == EXMEMALUOut[9:0] ? DMemory_243 : _GEN_1359; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1361 = 10'hf4 == EXMEMALUOut[9:0] ? DMemory_244 : _GEN_1360; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1362 = 10'hf5 == EXMEMALUOut[9:0] ? DMemory_245 : _GEN_1361; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1363 = 10'hf6 == EXMEMALUOut[9:0] ? DMemory_246 : _GEN_1362; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1364 = 10'hf7 == EXMEMALUOut[9:0] ? DMemory_247 : _GEN_1363; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1365 = 10'hf8 == EXMEMALUOut[9:0] ? DMemory_248 : _GEN_1364; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1366 = 10'hf9 == EXMEMALUOut[9:0] ? DMemory_249 : _GEN_1365; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1367 = 10'hfa == EXMEMALUOut[9:0] ? DMemory_250 : _GEN_1366; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1368 = 10'hfb == EXMEMALUOut[9:0] ? DMemory_251 : _GEN_1367; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1369 = 10'hfc == EXMEMALUOut[9:0] ? DMemory_252 : _GEN_1368; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1370 = 10'hfd == EXMEMALUOut[9:0] ? DMemory_253 : _GEN_1369; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1371 = 10'hfe == EXMEMALUOut[9:0] ? DMemory_254 : _GEN_1370; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1372 = 10'hff == EXMEMALUOut[9:0] ? DMemory_255 : _GEN_1371; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1373 = 10'h100 == EXMEMALUOut[9:0] ? DMemory_256 : _GEN_1372; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1374 = 10'h101 == EXMEMALUOut[9:0] ? DMemory_257 : _GEN_1373; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1375 = 10'h102 == EXMEMALUOut[9:0] ? DMemory_258 : _GEN_1374; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1376 = 10'h103 == EXMEMALUOut[9:0] ? DMemory_259 : _GEN_1375; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1377 = 10'h104 == EXMEMALUOut[9:0] ? DMemory_260 : _GEN_1376; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1378 = 10'h105 == EXMEMALUOut[9:0] ? DMemory_261 : _GEN_1377; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1379 = 10'h106 == EXMEMALUOut[9:0] ? DMemory_262 : _GEN_1378; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1380 = 10'h107 == EXMEMALUOut[9:0] ? DMemory_263 : _GEN_1379; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1381 = 10'h108 == EXMEMALUOut[9:0] ? DMemory_264 : _GEN_1380; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1382 = 10'h109 == EXMEMALUOut[9:0] ? DMemory_265 : _GEN_1381; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1383 = 10'h10a == EXMEMALUOut[9:0] ? DMemory_266 : _GEN_1382; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1384 = 10'h10b == EXMEMALUOut[9:0] ? DMemory_267 : _GEN_1383; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1385 = 10'h10c == EXMEMALUOut[9:0] ? DMemory_268 : _GEN_1384; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1386 = 10'h10d == EXMEMALUOut[9:0] ? DMemory_269 : _GEN_1385; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1387 = 10'h10e == EXMEMALUOut[9:0] ? DMemory_270 : _GEN_1386; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1388 = 10'h10f == EXMEMALUOut[9:0] ? DMemory_271 : _GEN_1387; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1389 = 10'h110 == EXMEMALUOut[9:0] ? DMemory_272 : _GEN_1388; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1390 = 10'h111 == EXMEMALUOut[9:0] ? DMemory_273 : _GEN_1389; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1391 = 10'h112 == EXMEMALUOut[9:0] ? DMemory_274 : _GEN_1390; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1392 = 10'h113 == EXMEMALUOut[9:0] ? DMemory_275 : _GEN_1391; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1393 = 10'h114 == EXMEMALUOut[9:0] ? DMemory_276 : _GEN_1392; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1394 = 10'h115 == EXMEMALUOut[9:0] ? DMemory_277 : _GEN_1393; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1395 = 10'h116 == EXMEMALUOut[9:0] ? DMemory_278 : _GEN_1394; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1396 = 10'h117 == EXMEMALUOut[9:0] ? DMemory_279 : _GEN_1395; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1397 = 10'h118 == EXMEMALUOut[9:0] ? DMemory_280 : _GEN_1396; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1398 = 10'h119 == EXMEMALUOut[9:0] ? DMemory_281 : _GEN_1397; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1399 = 10'h11a == EXMEMALUOut[9:0] ? DMemory_282 : _GEN_1398; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1400 = 10'h11b == EXMEMALUOut[9:0] ? DMemory_283 : _GEN_1399; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1401 = 10'h11c == EXMEMALUOut[9:0] ? DMemory_284 : _GEN_1400; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1402 = 10'h11d == EXMEMALUOut[9:0] ? DMemory_285 : _GEN_1401; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1403 = 10'h11e == EXMEMALUOut[9:0] ? DMemory_286 : _GEN_1402; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1404 = 10'h11f == EXMEMALUOut[9:0] ? DMemory_287 : _GEN_1403; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1405 = 10'h120 == EXMEMALUOut[9:0] ? DMemory_288 : _GEN_1404; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1406 = 10'h121 == EXMEMALUOut[9:0] ? DMemory_289 : _GEN_1405; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1407 = 10'h122 == EXMEMALUOut[9:0] ? DMemory_290 : _GEN_1406; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1408 = 10'h123 == EXMEMALUOut[9:0] ? DMemory_291 : _GEN_1407; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1409 = 10'h124 == EXMEMALUOut[9:0] ? DMemory_292 : _GEN_1408; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1410 = 10'h125 == EXMEMALUOut[9:0] ? DMemory_293 : _GEN_1409; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1411 = 10'h126 == EXMEMALUOut[9:0] ? DMemory_294 : _GEN_1410; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1412 = 10'h127 == EXMEMALUOut[9:0] ? DMemory_295 : _GEN_1411; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1413 = 10'h128 == EXMEMALUOut[9:0] ? DMemory_296 : _GEN_1412; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1414 = 10'h129 == EXMEMALUOut[9:0] ? DMemory_297 : _GEN_1413; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1415 = 10'h12a == EXMEMALUOut[9:0] ? DMemory_298 : _GEN_1414; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1416 = 10'h12b == EXMEMALUOut[9:0] ? DMemory_299 : _GEN_1415; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1417 = 10'h12c == EXMEMALUOut[9:0] ? DMemory_300 : _GEN_1416; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1418 = 10'h12d == EXMEMALUOut[9:0] ? DMemory_301 : _GEN_1417; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1419 = 10'h12e == EXMEMALUOut[9:0] ? DMemory_302 : _GEN_1418; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1420 = 10'h12f == EXMEMALUOut[9:0] ? DMemory_303 : _GEN_1419; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1421 = 10'h130 == EXMEMALUOut[9:0] ? DMemory_304 : _GEN_1420; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1422 = 10'h131 == EXMEMALUOut[9:0] ? DMemory_305 : _GEN_1421; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1423 = 10'h132 == EXMEMALUOut[9:0] ? DMemory_306 : _GEN_1422; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1424 = 10'h133 == EXMEMALUOut[9:0] ? DMemory_307 : _GEN_1423; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1425 = 10'h134 == EXMEMALUOut[9:0] ? DMemory_308 : _GEN_1424; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1426 = 10'h135 == EXMEMALUOut[9:0] ? DMemory_309 : _GEN_1425; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1427 = 10'h136 == EXMEMALUOut[9:0] ? DMemory_310 : _GEN_1426; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1428 = 10'h137 == EXMEMALUOut[9:0] ? DMemory_311 : _GEN_1427; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1429 = 10'h138 == EXMEMALUOut[9:0] ? DMemory_312 : _GEN_1428; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1430 = 10'h139 == EXMEMALUOut[9:0] ? DMemory_313 : _GEN_1429; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1431 = 10'h13a == EXMEMALUOut[9:0] ? DMemory_314 : _GEN_1430; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1432 = 10'h13b == EXMEMALUOut[9:0] ? DMemory_315 : _GEN_1431; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1433 = 10'h13c == EXMEMALUOut[9:0] ? DMemory_316 : _GEN_1432; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1434 = 10'h13d == EXMEMALUOut[9:0] ? DMemory_317 : _GEN_1433; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1435 = 10'h13e == EXMEMALUOut[9:0] ? DMemory_318 : _GEN_1434; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1436 = 10'h13f == EXMEMALUOut[9:0] ? DMemory_319 : _GEN_1435; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1437 = 10'h140 == EXMEMALUOut[9:0] ? DMemory_320 : _GEN_1436; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1438 = 10'h141 == EXMEMALUOut[9:0] ? DMemory_321 : _GEN_1437; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1439 = 10'h142 == EXMEMALUOut[9:0] ? DMemory_322 : _GEN_1438; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1440 = 10'h143 == EXMEMALUOut[9:0] ? DMemory_323 : _GEN_1439; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1441 = 10'h144 == EXMEMALUOut[9:0] ? DMemory_324 : _GEN_1440; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1442 = 10'h145 == EXMEMALUOut[9:0] ? DMemory_325 : _GEN_1441; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1443 = 10'h146 == EXMEMALUOut[9:0] ? DMemory_326 : _GEN_1442; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1444 = 10'h147 == EXMEMALUOut[9:0] ? DMemory_327 : _GEN_1443; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1445 = 10'h148 == EXMEMALUOut[9:0] ? DMemory_328 : _GEN_1444; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1446 = 10'h149 == EXMEMALUOut[9:0] ? DMemory_329 : _GEN_1445; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1447 = 10'h14a == EXMEMALUOut[9:0] ? DMemory_330 : _GEN_1446; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1448 = 10'h14b == EXMEMALUOut[9:0] ? DMemory_331 : _GEN_1447; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1449 = 10'h14c == EXMEMALUOut[9:0] ? DMemory_332 : _GEN_1448; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1450 = 10'h14d == EXMEMALUOut[9:0] ? DMemory_333 : _GEN_1449; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1451 = 10'h14e == EXMEMALUOut[9:0] ? DMemory_334 : _GEN_1450; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1452 = 10'h14f == EXMEMALUOut[9:0] ? DMemory_335 : _GEN_1451; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1453 = 10'h150 == EXMEMALUOut[9:0] ? DMemory_336 : _GEN_1452; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1454 = 10'h151 == EXMEMALUOut[9:0] ? DMemory_337 : _GEN_1453; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1455 = 10'h152 == EXMEMALUOut[9:0] ? DMemory_338 : _GEN_1454; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1456 = 10'h153 == EXMEMALUOut[9:0] ? DMemory_339 : _GEN_1455; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1457 = 10'h154 == EXMEMALUOut[9:0] ? DMemory_340 : _GEN_1456; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1458 = 10'h155 == EXMEMALUOut[9:0] ? DMemory_341 : _GEN_1457; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1459 = 10'h156 == EXMEMALUOut[9:0] ? DMemory_342 : _GEN_1458; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1460 = 10'h157 == EXMEMALUOut[9:0] ? DMemory_343 : _GEN_1459; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1461 = 10'h158 == EXMEMALUOut[9:0] ? DMemory_344 : _GEN_1460; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1462 = 10'h159 == EXMEMALUOut[9:0] ? DMemory_345 : _GEN_1461; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1463 = 10'h15a == EXMEMALUOut[9:0] ? DMemory_346 : _GEN_1462; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1464 = 10'h15b == EXMEMALUOut[9:0] ? DMemory_347 : _GEN_1463; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1465 = 10'h15c == EXMEMALUOut[9:0] ? DMemory_348 : _GEN_1464; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1466 = 10'h15d == EXMEMALUOut[9:0] ? DMemory_349 : _GEN_1465; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1467 = 10'h15e == EXMEMALUOut[9:0] ? DMemory_350 : _GEN_1466; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1468 = 10'h15f == EXMEMALUOut[9:0] ? DMemory_351 : _GEN_1467; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1469 = 10'h160 == EXMEMALUOut[9:0] ? DMemory_352 : _GEN_1468; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1470 = 10'h161 == EXMEMALUOut[9:0] ? DMemory_353 : _GEN_1469; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1471 = 10'h162 == EXMEMALUOut[9:0] ? DMemory_354 : _GEN_1470; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1472 = 10'h163 == EXMEMALUOut[9:0] ? DMemory_355 : _GEN_1471; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1473 = 10'h164 == EXMEMALUOut[9:0] ? DMemory_356 : _GEN_1472; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1474 = 10'h165 == EXMEMALUOut[9:0] ? DMemory_357 : _GEN_1473; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1475 = 10'h166 == EXMEMALUOut[9:0] ? DMemory_358 : _GEN_1474; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1476 = 10'h167 == EXMEMALUOut[9:0] ? DMemory_359 : _GEN_1475; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1477 = 10'h168 == EXMEMALUOut[9:0] ? DMemory_360 : _GEN_1476; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1478 = 10'h169 == EXMEMALUOut[9:0] ? DMemory_361 : _GEN_1477; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1479 = 10'h16a == EXMEMALUOut[9:0] ? DMemory_362 : _GEN_1478; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1480 = 10'h16b == EXMEMALUOut[9:0] ? DMemory_363 : _GEN_1479; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1481 = 10'h16c == EXMEMALUOut[9:0] ? DMemory_364 : _GEN_1480; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1482 = 10'h16d == EXMEMALUOut[9:0] ? DMemory_365 : _GEN_1481; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1483 = 10'h16e == EXMEMALUOut[9:0] ? DMemory_366 : _GEN_1482; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1484 = 10'h16f == EXMEMALUOut[9:0] ? DMemory_367 : _GEN_1483; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1485 = 10'h170 == EXMEMALUOut[9:0] ? DMemory_368 : _GEN_1484; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1486 = 10'h171 == EXMEMALUOut[9:0] ? DMemory_369 : _GEN_1485; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1487 = 10'h172 == EXMEMALUOut[9:0] ? DMemory_370 : _GEN_1486; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1488 = 10'h173 == EXMEMALUOut[9:0] ? DMemory_371 : _GEN_1487; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1489 = 10'h174 == EXMEMALUOut[9:0] ? DMemory_372 : _GEN_1488; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1490 = 10'h175 == EXMEMALUOut[9:0] ? DMemory_373 : _GEN_1489; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1491 = 10'h176 == EXMEMALUOut[9:0] ? DMemory_374 : _GEN_1490; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1492 = 10'h177 == EXMEMALUOut[9:0] ? DMemory_375 : _GEN_1491; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1493 = 10'h178 == EXMEMALUOut[9:0] ? DMemory_376 : _GEN_1492; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1494 = 10'h179 == EXMEMALUOut[9:0] ? DMemory_377 : _GEN_1493; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1495 = 10'h17a == EXMEMALUOut[9:0] ? DMemory_378 : _GEN_1494; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1496 = 10'h17b == EXMEMALUOut[9:0] ? DMemory_379 : _GEN_1495; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1497 = 10'h17c == EXMEMALUOut[9:0] ? DMemory_380 : _GEN_1496; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1498 = 10'h17d == EXMEMALUOut[9:0] ? DMemory_381 : _GEN_1497; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1499 = 10'h17e == EXMEMALUOut[9:0] ? DMemory_382 : _GEN_1498; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1500 = 10'h17f == EXMEMALUOut[9:0] ? DMemory_383 : _GEN_1499; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1501 = 10'h180 == EXMEMALUOut[9:0] ? DMemory_384 : _GEN_1500; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1502 = 10'h181 == EXMEMALUOut[9:0] ? DMemory_385 : _GEN_1501; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1503 = 10'h182 == EXMEMALUOut[9:0] ? DMemory_386 : _GEN_1502; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1504 = 10'h183 == EXMEMALUOut[9:0] ? DMemory_387 : _GEN_1503; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1505 = 10'h184 == EXMEMALUOut[9:0] ? DMemory_388 : _GEN_1504; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1506 = 10'h185 == EXMEMALUOut[9:0] ? DMemory_389 : _GEN_1505; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1507 = 10'h186 == EXMEMALUOut[9:0] ? DMemory_390 : _GEN_1506; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1508 = 10'h187 == EXMEMALUOut[9:0] ? DMemory_391 : _GEN_1507; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1509 = 10'h188 == EXMEMALUOut[9:0] ? DMemory_392 : _GEN_1508; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1510 = 10'h189 == EXMEMALUOut[9:0] ? DMemory_393 : _GEN_1509; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1511 = 10'h18a == EXMEMALUOut[9:0] ? DMemory_394 : _GEN_1510; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1512 = 10'h18b == EXMEMALUOut[9:0] ? DMemory_395 : _GEN_1511; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1513 = 10'h18c == EXMEMALUOut[9:0] ? DMemory_396 : _GEN_1512; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1514 = 10'h18d == EXMEMALUOut[9:0] ? DMemory_397 : _GEN_1513; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1515 = 10'h18e == EXMEMALUOut[9:0] ? DMemory_398 : _GEN_1514; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1516 = 10'h18f == EXMEMALUOut[9:0] ? DMemory_399 : _GEN_1515; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1517 = 10'h190 == EXMEMALUOut[9:0] ? DMemory_400 : _GEN_1516; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1518 = 10'h191 == EXMEMALUOut[9:0] ? DMemory_401 : _GEN_1517; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1519 = 10'h192 == EXMEMALUOut[9:0] ? DMemory_402 : _GEN_1518; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1520 = 10'h193 == EXMEMALUOut[9:0] ? DMemory_403 : _GEN_1519; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1521 = 10'h194 == EXMEMALUOut[9:0] ? DMemory_404 : _GEN_1520; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1522 = 10'h195 == EXMEMALUOut[9:0] ? DMemory_405 : _GEN_1521; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1523 = 10'h196 == EXMEMALUOut[9:0] ? DMemory_406 : _GEN_1522; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1524 = 10'h197 == EXMEMALUOut[9:0] ? DMemory_407 : _GEN_1523; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1525 = 10'h198 == EXMEMALUOut[9:0] ? DMemory_408 : _GEN_1524; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1526 = 10'h199 == EXMEMALUOut[9:0] ? DMemory_409 : _GEN_1525; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1527 = 10'h19a == EXMEMALUOut[9:0] ? DMemory_410 : _GEN_1526; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1528 = 10'h19b == EXMEMALUOut[9:0] ? DMemory_411 : _GEN_1527; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1529 = 10'h19c == EXMEMALUOut[9:0] ? DMemory_412 : _GEN_1528; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1530 = 10'h19d == EXMEMALUOut[9:0] ? DMemory_413 : _GEN_1529; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1531 = 10'h19e == EXMEMALUOut[9:0] ? DMemory_414 : _GEN_1530; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1532 = 10'h19f == EXMEMALUOut[9:0] ? DMemory_415 : _GEN_1531; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1533 = 10'h1a0 == EXMEMALUOut[9:0] ? DMemory_416 : _GEN_1532; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1534 = 10'h1a1 == EXMEMALUOut[9:0] ? DMemory_417 : _GEN_1533; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1535 = 10'h1a2 == EXMEMALUOut[9:0] ? DMemory_418 : _GEN_1534; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1536 = 10'h1a3 == EXMEMALUOut[9:0] ? DMemory_419 : _GEN_1535; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1537 = 10'h1a4 == EXMEMALUOut[9:0] ? DMemory_420 : _GEN_1536; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1538 = 10'h1a5 == EXMEMALUOut[9:0] ? DMemory_421 : _GEN_1537; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1539 = 10'h1a6 == EXMEMALUOut[9:0] ? DMemory_422 : _GEN_1538; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1540 = 10'h1a7 == EXMEMALUOut[9:0] ? DMemory_423 : _GEN_1539; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1541 = 10'h1a8 == EXMEMALUOut[9:0] ? DMemory_424 : _GEN_1540; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1542 = 10'h1a9 == EXMEMALUOut[9:0] ? DMemory_425 : _GEN_1541; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1543 = 10'h1aa == EXMEMALUOut[9:0] ? DMemory_426 : _GEN_1542; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1544 = 10'h1ab == EXMEMALUOut[9:0] ? DMemory_427 : _GEN_1543; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1545 = 10'h1ac == EXMEMALUOut[9:0] ? DMemory_428 : _GEN_1544; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1546 = 10'h1ad == EXMEMALUOut[9:0] ? DMemory_429 : _GEN_1545; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1547 = 10'h1ae == EXMEMALUOut[9:0] ? DMemory_430 : _GEN_1546; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1548 = 10'h1af == EXMEMALUOut[9:0] ? DMemory_431 : _GEN_1547; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1549 = 10'h1b0 == EXMEMALUOut[9:0] ? DMemory_432 : _GEN_1548; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1550 = 10'h1b1 == EXMEMALUOut[9:0] ? DMemory_433 : _GEN_1549; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1551 = 10'h1b2 == EXMEMALUOut[9:0] ? DMemory_434 : _GEN_1550; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1552 = 10'h1b3 == EXMEMALUOut[9:0] ? DMemory_435 : _GEN_1551; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1553 = 10'h1b4 == EXMEMALUOut[9:0] ? DMemory_436 : _GEN_1552; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1554 = 10'h1b5 == EXMEMALUOut[9:0] ? DMemory_437 : _GEN_1553; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1555 = 10'h1b6 == EXMEMALUOut[9:0] ? DMemory_438 : _GEN_1554; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1556 = 10'h1b7 == EXMEMALUOut[9:0] ? DMemory_439 : _GEN_1555; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1557 = 10'h1b8 == EXMEMALUOut[9:0] ? DMemory_440 : _GEN_1556; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1558 = 10'h1b9 == EXMEMALUOut[9:0] ? DMemory_441 : _GEN_1557; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1559 = 10'h1ba == EXMEMALUOut[9:0] ? DMemory_442 : _GEN_1558; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1560 = 10'h1bb == EXMEMALUOut[9:0] ? DMemory_443 : _GEN_1559; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1561 = 10'h1bc == EXMEMALUOut[9:0] ? DMemory_444 : _GEN_1560; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1562 = 10'h1bd == EXMEMALUOut[9:0] ? DMemory_445 : _GEN_1561; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1563 = 10'h1be == EXMEMALUOut[9:0] ? DMemory_446 : _GEN_1562; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1564 = 10'h1bf == EXMEMALUOut[9:0] ? DMemory_447 : _GEN_1563; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1565 = 10'h1c0 == EXMEMALUOut[9:0] ? DMemory_448 : _GEN_1564; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1566 = 10'h1c1 == EXMEMALUOut[9:0] ? DMemory_449 : _GEN_1565; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1567 = 10'h1c2 == EXMEMALUOut[9:0] ? DMemory_450 : _GEN_1566; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1568 = 10'h1c3 == EXMEMALUOut[9:0] ? DMemory_451 : _GEN_1567; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1569 = 10'h1c4 == EXMEMALUOut[9:0] ? DMemory_452 : _GEN_1568; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1570 = 10'h1c5 == EXMEMALUOut[9:0] ? DMemory_453 : _GEN_1569; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1571 = 10'h1c6 == EXMEMALUOut[9:0] ? DMemory_454 : _GEN_1570; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1572 = 10'h1c7 == EXMEMALUOut[9:0] ? DMemory_455 : _GEN_1571; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1573 = 10'h1c8 == EXMEMALUOut[9:0] ? DMemory_456 : _GEN_1572; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1574 = 10'h1c9 == EXMEMALUOut[9:0] ? DMemory_457 : _GEN_1573; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1575 = 10'h1ca == EXMEMALUOut[9:0] ? DMemory_458 : _GEN_1574; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1576 = 10'h1cb == EXMEMALUOut[9:0] ? DMemory_459 : _GEN_1575; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1577 = 10'h1cc == EXMEMALUOut[9:0] ? DMemory_460 : _GEN_1576; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1578 = 10'h1cd == EXMEMALUOut[9:0] ? DMemory_461 : _GEN_1577; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1579 = 10'h1ce == EXMEMALUOut[9:0] ? DMemory_462 : _GEN_1578; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1580 = 10'h1cf == EXMEMALUOut[9:0] ? DMemory_463 : _GEN_1579; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1581 = 10'h1d0 == EXMEMALUOut[9:0] ? DMemory_464 : _GEN_1580; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1582 = 10'h1d1 == EXMEMALUOut[9:0] ? DMemory_465 : _GEN_1581; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1583 = 10'h1d2 == EXMEMALUOut[9:0] ? DMemory_466 : _GEN_1582; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1584 = 10'h1d3 == EXMEMALUOut[9:0] ? DMemory_467 : _GEN_1583; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1585 = 10'h1d4 == EXMEMALUOut[9:0] ? DMemory_468 : _GEN_1584; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1586 = 10'h1d5 == EXMEMALUOut[9:0] ? DMemory_469 : _GEN_1585; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1587 = 10'h1d6 == EXMEMALUOut[9:0] ? DMemory_470 : _GEN_1586; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1588 = 10'h1d7 == EXMEMALUOut[9:0] ? DMemory_471 : _GEN_1587; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1589 = 10'h1d8 == EXMEMALUOut[9:0] ? DMemory_472 : _GEN_1588; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1590 = 10'h1d9 == EXMEMALUOut[9:0] ? DMemory_473 : _GEN_1589; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1591 = 10'h1da == EXMEMALUOut[9:0] ? DMemory_474 : _GEN_1590; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1592 = 10'h1db == EXMEMALUOut[9:0] ? DMemory_475 : _GEN_1591; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1593 = 10'h1dc == EXMEMALUOut[9:0] ? DMemory_476 : _GEN_1592; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1594 = 10'h1dd == EXMEMALUOut[9:0] ? DMemory_477 : _GEN_1593; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1595 = 10'h1de == EXMEMALUOut[9:0] ? DMemory_478 : _GEN_1594; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1596 = 10'h1df == EXMEMALUOut[9:0] ? DMemory_479 : _GEN_1595; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1597 = 10'h1e0 == EXMEMALUOut[9:0] ? DMemory_480 : _GEN_1596; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1598 = 10'h1e1 == EXMEMALUOut[9:0] ? DMemory_481 : _GEN_1597; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1599 = 10'h1e2 == EXMEMALUOut[9:0] ? DMemory_482 : _GEN_1598; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1600 = 10'h1e3 == EXMEMALUOut[9:0] ? DMemory_483 : _GEN_1599; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1601 = 10'h1e4 == EXMEMALUOut[9:0] ? DMemory_484 : _GEN_1600; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1602 = 10'h1e5 == EXMEMALUOut[9:0] ? DMemory_485 : _GEN_1601; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1603 = 10'h1e6 == EXMEMALUOut[9:0] ? DMemory_486 : _GEN_1602; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1604 = 10'h1e7 == EXMEMALUOut[9:0] ? DMemory_487 : _GEN_1603; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1605 = 10'h1e8 == EXMEMALUOut[9:0] ? DMemory_488 : _GEN_1604; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1606 = 10'h1e9 == EXMEMALUOut[9:0] ? DMemory_489 : _GEN_1605; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1607 = 10'h1ea == EXMEMALUOut[9:0] ? DMemory_490 : _GEN_1606; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1608 = 10'h1eb == EXMEMALUOut[9:0] ? DMemory_491 : _GEN_1607; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1609 = 10'h1ec == EXMEMALUOut[9:0] ? DMemory_492 : _GEN_1608; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1610 = 10'h1ed == EXMEMALUOut[9:0] ? DMemory_493 : _GEN_1609; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1611 = 10'h1ee == EXMEMALUOut[9:0] ? DMemory_494 : _GEN_1610; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1612 = 10'h1ef == EXMEMALUOut[9:0] ? DMemory_495 : _GEN_1611; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1613 = 10'h1f0 == EXMEMALUOut[9:0] ? DMemory_496 : _GEN_1612; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1614 = 10'h1f1 == EXMEMALUOut[9:0] ? DMemory_497 : _GEN_1613; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1615 = 10'h1f2 == EXMEMALUOut[9:0] ? DMemory_498 : _GEN_1614; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1616 = 10'h1f3 == EXMEMALUOut[9:0] ? DMemory_499 : _GEN_1615; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1617 = 10'h1f4 == EXMEMALUOut[9:0] ? DMemory_500 : _GEN_1616; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1618 = 10'h1f5 == EXMEMALUOut[9:0] ? DMemory_501 : _GEN_1617; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1619 = 10'h1f6 == EXMEMALUOut[9:0] ? DMemory_502 : _GEN_1618; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1620 = 10'h1f7 == EXMEMALUOut[9:0] ? DMemory_503 : _GEN_1619; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1621 = 10'h1f8 == EXMEMALUOut[9:0] ? DMemory_504 : _GEN_1620; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1622 = 10'h1f9 == EXMEMALUOut[9:0] ? DMemory_505 : _GEN_1621; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1623 = 10'h1fa == EXMEMALUOut[9:0] ? DMemory_506 : _GEN_1622; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1624 = 10'h1fb == EXMEMALUOut[9:0] ? DMemory_507 : _GEN_1623; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1625 = 10'h1fc == EXMEMALUOut[9:0] ? DMemory_508 : _GEN_1624; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1626 = 10'h1fd == EXMEMALUOut[9:0] ? DMemory_509 : _GEN_1625; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1627 = 10'h1fe == EXMEMALUOut[9:0] ? DMemory_510 : _GEN_1626; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1628 = 10'h1ff == EXMEMALUOut[9:0] ? DMemory_511 : _GEN_1627; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1629 = 10'h200 == EXMEMALUOut[9:0] ? DMemory_512 : _GEN_1628; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1630 = 10'h201 == EXMEMALUOut[9:0] ? DMemory_513 : _GEN_1629; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1631 = 10'h202 == EXMEMALUOut[9:0] ? DMemory_514 : _GEN_1630; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1632 = 10'h203 == EXMEMALUOut[9:0] ? DMemory_515 : _GEN_1631; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1633 = 10'h204 == EXMEMALUOut[9:0] ? DMemory_516 : _GEN_1632; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1634 = 10'h205 == EXMEMALUOut[9:0] ? DMemory_517 : _GEN_1633; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1635 = 10'h206 == EXMEMALUOut[9:0] ? DMemory_518 : _GEN_1634; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1636 = 10'h207 == EXMEMALUOut[9:0] ? DMemory_519 : _GEN_1635; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1637 = 10'h208 == EXMEMALUOut[9:0] ? DMemory_520 : _GEN_1636; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1638 = 10'h209 == EXMEMALUOut[9:0] ? DMemory_521 : _GEN_1637; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1639 = 10'h20a == EXMEMALUOut[9:0] ? DMemory_522 : _GEN_1638; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1640 = 10'h20b == EXMEMALUOut[9:0] ? DMemory_523 : _GEN_1639; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1641 = 10'h20c == EXMEMALUOut[9:0] ? DMemory_524 : _GEN_1640; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1642 = 10'h20d == EXMEMALUOut[9:0] ? DMemory_525 : _GEN_1641; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1643 = 10'h20e == EXMEMALUOut[9:0] ? DMemory_526 : _GEN_1642; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1644 = 10'h20f == EXMEMALUOut[9:0] ? DMemory_527 : _GEN_1643; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1645 = 10'h210 == EXMEMALUOut[9:0] ? DMemory_528 : _GEN_1644; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1646 = 10'h211 == EXMEMALUOut[9:0] ? DMemory_529 : _GEN_1645; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1647 = 10'h212 == EXMEMALUOut[9:0] ? DMemory_530 : _GEN_1646; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1648 = 10'h213 == EXMEMALUOut[9:0] ? DMemory_531 : _GEN_1647; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1649 = 10'h214 == EXMEMALUOut[9:0] ? DMemory_532 : _GEN_1648; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1650 = 10'h215 == EXMEMALUOut[9:0] ? DMemory_533 : _GEN_1649; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1651 = 10'h216 == EXMEMALUOut[9:0] ? DMemory_534 : _GEN_1650; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1652 = 10'h217 == EXMEMALUOut[9:0] ? DMemory_535 : _GEN_1651; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1653 = 10'h218 == EXMEMALUOut[9:0] ? DMemory_536 : _GEN_1652; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1654 = 10'h219 == EXMEMALUOut[9:0] ? DMemory_537 : _GEN_1653; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1655 = 10'h21a == EXMEMALUOut[9:0] ? DMemory_538 : _GEN_1654; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1656 = 10'h21b == EXMEMALUOut[9:0] ? DMemory_539 : _GEN_1655; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1657 = 10'h21c == EXMEMALUOut[9:0] ? DMemory_540 : _GEN_1656; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1658 = 10'h21d == EXMEMALUOut[9:0] ? DMemory_541 : _GEN_1657; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1659 = 10'h21e == EXMEMALUOut[9:0] ? DMemory_542 : _GEN_1658; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1660 = 10'h21f == EXMEMALUOut[9:0] ? DMemory_543 : _GEN_1659; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1661 = 10'h220 == EXMEMALUOut[9:0] ? DMemory_544 : _GEN_1660; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1662 = 10'h221 == EXMEMALUOut[9:0] ? DMemory_545 : _GEN_1661; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1663 = 10'h222 == EXMEMALUOut[9:0] ? DMemory_546 : _GEN_1662; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1664 = 10'h223 == EXMEMALUOut[9:0] ? DMemory_547 : _GEN_1663; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1665 = 10'h224 == EXMEMALUOut[9:0] ? DMemory_548 : _GEN_1664; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1666 = 10'h225 == EXMEMALUOut[9:0] ? DMemory_549 : _GEN_1665; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1667 = 10'h226 == EXMEMALUOut[9:0] ? DMemory_550 : _GEN_1666; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1668 = 10'h227 == EXMEMALUOut[9:0] ? DMemory_551 : _GEN_1667; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1669 = 10'h228 == EXMEMALUOut[9:0] ? DMemory_552 : _GEN_1668; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1670 = 10'h229 == EXMEMALUOut[9:0] ? DMemory_553 : _GEN_1669; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1671 = 10'h22a == EXMEMALUOut[9:0] ? DMemory_554 : _GEN_1670; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1672 = 10'h22b == EXMEMALUOut[9:0] ? DMemory_555 : _GEN_1671; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1673 = 10'h22c == EXMEMALUOut[9:0] ? DMemory_556 : _GEN_1672; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1674 = 10'h22d == EXMEMALUOut[9:0] ? DMemory_557 : _GEN_1673; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1675 = 10'h22e == EXMEMALUOut[9:0] ? DMemory_558 : _GEN_1674; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1676 = 10'h22f == EXMEMALUOut[9:0] ? DMemory_559 : _GEN_1675; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1677 = 10'h230 == EXMEMALUOut[9:0] ? DMemory_560 : _GEN_1676; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1678 = 10'h231 == EXMEMALUOut[9:0] ? DMemory_561 : _GEN_1677; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1679 = 10'h232 == EXMEMALUOut[9:0] ? DMemory_562 : _GEN_1678; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1680 = 10'h233 == EXMEMALUOut[9:0] ? DMemory_563 : _GEN_1679; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1681 = 10'h234 == EXMEMALUOut[9:0] ? DMemory_564 : _GEN_1680; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1682 = 10'h235 == EXMEMALUOut[9:0] ? DMemory_565 : _GEN_1681; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1683 = 10'h236 == EXMEMALUOut[9:0] ? DMemory_566 : _GEN_1682; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1684 = 10'h237 == EXMEMALUOut[9:0] ? DMemory_567 : _GEN_1683; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1685 = 10'h238 == EXMEMALUOut[9:0] ? DMemory_568 : _GEN_1684; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1686 = 10'h239 == EXMEMALUOut[9:0] ? DMemory_569 : _GEN_1685; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1687 = 10'h23a == EXMEMALUOut[9:0] ? DMemory_570 : _GEN_1686; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1688 = 10'h23b == EXMEMALUOut[9:0] ? DMemory_571 : _GEN_1687; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1689 = 10'h23c == EXMEMALUOut[9:0] ? DMemory_572 : _GEN_1688; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1690 = 10'h23d == EXMEMALUOut[9:0] ? DMemory_573 : _GEN_1689; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1691 = 10'h23e == EXMEMALUOut[9:0] ? DMemory_574 : _GEN_1690; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1692 = 10'h23f == EXMEMALUOut[9:0] ? DMemory_575 : _GEN_1691; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1693 = 10'h240 == EXMEMALUOut[9:0] ? DMemory_576 : _GEN_1692; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1694 = 10'h241 == EXMEMALUOut[9:0] ? DMemory_577 : _GEN_1693; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1695 = 10'h242 == EXMEMALUOut[9:0] ? DMemory_578 : _GEN_1694; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1696 = 10'h243 == EXMEMALUOut[9:0] ? DMemory_579 : _GEN_1695; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1697 = 10'h244 == EXMEMALUOut[9:0] ? DMemory_580 : _GEN_1696; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1698 = 10'h245 == EXMEMALUOut[9:0] ? DMemory_581 : _GEN_1697; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1699 = 10'h246 == EXMEMALUOut[9:0] ? DMemory_582 : _GEN_1698; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1700 = 10'h247 == EXMEMALUOut[9:0] ? DMemory_583 : _GEN_1699; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1701 = 10'h248 == EXMEMALUOut[9:0] ? DMemory_584 : _GEN_1700; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1702 = 10'h249 == EXMEMALUOut[9:0] ? DMemory_585 : _GEN_1701; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1703 = 10'h24a == EXMEMALUOut[9:0] ? DMemory_586 : _GEN_1702; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1704 = 10'h24b == EXMEMALUOut[9:0] ? DMemory_587 : _GEN_1703; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1705 = 10'h24c == EXMEMALUOut[9:0] ? DMemory_588 : _GEN_1704; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1706 = 10'h24d == EXMEMALUOut[9:0] ? DMemory_589 : _GEN_1705; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1707 = 10'h24e == EXMEMALUOut[9:0] ? DMemory_590 : _GEN_1706; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1708 = 10'h24f == EXMEMALUOut[9:0] ? DMemory_591 : _GEN_1707; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1709 = 10'h250 == EXMEMALUOut[9:0] ? DMemory_592 : _GEN_1708; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1710 = 10'h251 == EXMEMALUOut[9:0] ? DMemory_593 : _GEN_1709; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1711 = 10'h252 == EXMEMALUOut[9:0] ? DMemory_594 : _GEN_1710; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1712 = 10'h253 == EXMEMALUOut[9:0] ? DMemory_595 : _GEN_1711; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1713 = 10'h254 == EXMEMALUOut[9:0] ? DMemory_596 : _GEN_1712; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1714 = 10'h255 == EXMEMALUOut[9:0] ? DMemory_597 : _GEN_1713; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1715 = 10'h256 == EXMEMALUOut[9:0] ? DMemory_598 : _GEN_1714; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1716 = 10'h257 == EXMEMALUOut[9:0] ? DMemory_599 : _GEN_1715; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1717 = 10'h258 == EXMEMALUOut[9:0] ? DMemory_600 : _GEN_1716; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1718 = 10'h259 == EXMEMALUOut[9:0] ? DMemory_601 : _GEN_1717; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1719 = 10'h25a == EXMEMALUOut[9:0] ? DMemory_602 : _GEN_1718; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1720 = 10'h25b == EXMEMALUOut[9:0] ? DMemory_603 : _GEN_1719; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1721 = 10'h25c == EXMEMALUOut[9:0] ? DMemory_604 : _GEN_1720; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1722 = 10'h25d == EXMEMALUOut[9:0] ? DMemory_605 : _GEN_1721; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1723 = 10'h25e == EXMEMALUOut[9:0] ? DMemory_606 : _GEN_1722; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1724 = 10'h25f == EXMEMALUOut[9:0] ? DMemory_607 : _GEN_1723; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1725 = 10'h260 == EXMEMALUOut[9:0] ? DMemory_608 : _GEN_1724; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1726 = 10'h261 == EXMEMALUOut[9:0] ? DMemory_609 : _GEN_1725; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1727 = 10'h262 == EXMEMALUOut[9:0] ? DMemory_610 : _GEN_1726; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1728 = 10'h263 == EXMEMALUOut[9:0] ? DMemory_611 : _GEN_1727; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1729 = 10'h264 == EXMEMALUOut[9:0] ? DMemory_612 : _GEN_1728; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1730 = 10'h265 == EXMEMALUOut[9:0] ? DMemory_613 : _GEN_1729; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1731 = 10'h266 == EXMEMALUOut[9:0] ? DMemory_614 : _GEN_1730; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1732 = 10'h267 == EXMEMALUOut[9:0] ? DMemory_615 : _GEN_1731; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1733 = 10'h268 == EXMEMALUOut[9:0] ? DMemory_616 : _GEN_1732; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1734 = 10'h269 == EXMEMALUOut[9:0] ? DMemory_617 : _GEN_1733; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1735 = 10'h26a == EXMEMALUOut[9:0] ? DMemory_618 : _GEN_1734; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1736 = 10'h26b == EXMEMALUOut[9:0] ? DMemory_619 : _GEN_1735; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1737 = 10'h26c == EXMEMALUOut[9:0] ? DMemory_620 : _GEN_1736; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1738 = 10'h26d == EXMEMALUOut[9:0] ? DMemory_621 : _GEN_1737; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1739 = 10'h26e == EXMEMALUOut[9:0] ? DMemory_622 : _GEN_1738; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1740 = 10'h26f == EXMEMALUOut[9:0] ? DMemory_623 : _GEN_1739; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1741 = 10'h270 == EXMEMALUOut[9:0] ? DMemory_624 : _GEN_1740; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1742 = 10'h271 == EXMEMALUOut[9:0] ? DMemory_625 : _GEN_1741; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1743 = 10'h272 == EXMEMALUOut[9:0] ? DMemory_626 : _GEN_1742; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1744 = 10'h273 == EXMEMALUOut[9:0] ? DMemory_627 : _GEN_1743; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1745 = 10'h274 == EXMEMALUOut[9:0] ? DMemory_628 : _GEN_1744; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1746 = 10'h275 == EXMEMALUOut[9:0] ? DMemory_629 : _GEN_1745; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1747 = 10'h276 == EXMEMALUOut[9:0] ? DMemory_630 : _GEN_1746; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1748 = 10'h277 == EXMEMALUOut[9:0] ? DMemory_631 : _GEN_1747; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1749 = 10'h278 == EXMEMALUOut[9:0] ? DMemory_632 : _GEN_1748; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1750 = 10'h279 == EXMEMALUOut[9:0] ? DMemory_633 : _GEN_1749; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1751 = 10'h27a == EXMEMALUOut[9:0] ? DMemory_634 : _GEN_1750; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1752 = 10'h27b == EXMEMALUOut[9:0] ? DMemory_635 : _GEN_1751; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1753 = 10'h27c == EXMEMALUOut[9:0] ? DMemory_636 : _GEN_1752; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1754 = 10'h27d == EXMEMALUOut[9:0] ? DMemory_637 : _GEN_1753; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1755 = 10'h27e == EXMEMALUOut[9:0] ? DMemory_638 : _GEN_1754; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1756 = 10'h27f == EXMEMALUOut[9:0] ? DMemory_639 : _GEN_1755; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1757 = 10'h280 == EXMEMALUOut[9:0] ? DMemory_640 : _GEN_1756; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1758 = 10'h281 == EXMEMALUOut[9:0] ? DMemory_641 : _GEN_1757; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1759 = 10'h282 == EXMEMALUOut[9:0] ? DMemory_642 : _GEN_1758; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1760 = 10'h283 == EXMEMALUOut[9:0] ? DMemory_643 : _GEN_1759; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1761 = 10'h284 == EXMEMALUOut[9:0] ? DMemory_644 : _GEN_1760; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1762 = 10'h285 == EXMEMALUOut[9:0] ? DMemory_645 : _GEN_1761; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1763 = 10'h286 == EXMEMALUOut[9:0] ? DMemory_646 : _GEN_1762; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1764 = 10'h287 == EXMEMALUOut[9:0] ? DMemory_647 : _GEN_1763; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1765 = 10'h288 == EXMEMALUOut[9:0] ? DMemory_648 : _GEN_1764; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1766 = 10'h289 == EXMEMALUOut[9:0] ? DMemory_649 : _GEN_1765; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1767 = 10'h28a == EXMEMALUOut[9:0] ? DMemory_650 : _GEN_1766; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1768 = 10'h28b == EXMEMALUOut[9:0] ? DMemory_651 : _GEN_1767; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1769 = 10'h28c == EXMEMALUOut[9:0] ? DMemory_652 : _GEN_1768; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1770 = 10'h28d == EXMEMALUOut[9:0] ? DMemory_653 : _GEN_1769; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1771 = 10'h28e == EXMEMALUOut[9:0] ? DMemory_654 : _GEN_1770; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1772 = 10'h28f == EXMEMALUOut[9:0] ? DMemory_655 : _GEN_1771; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1773 = 10'h290 == EXMEMALUOut[9:0] ? DMemory_656 : _GEN_1772; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1774 = 10'h291 == EXMEMALUOut[9:0] ? DMemory_657 : _GEN_1773; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1775 = 10'h292 == EXMEMALUOut[9:0] ? DMemory_658 : _GEN_1774; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1776 = 10'h293 == EXMEMALUOut[9:0] ? DMemory_659 : _GEN_1775; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1777 = 10'h294 == EXMEMALUOut[9:0] ? DMemory_660 : _GEN_1776; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1778 = 10'h295 == EXMEMALUOut[9:0] ? DMemory_661 : _GEN_1777; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1779 = 10'h296 == EXMEMALUOut[9:0] ? DMemory_662 : _GEN_1778; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1780 = 10'h297 == EXMEMALUOut[9:0] ? DMemory_663 : _GEN_1779; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1781 = 10'h298 == EXMEMALUOut[9:0] ? DMemory_664 : _GEN_1780; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1782 = 10'h299 == EXMEMALUOut[9:0] ? DMemory_665 : _GEN_1781; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1783 = 10'h29a == EXMEMALUOut[9:0] ? DMemory_666 : _GEN_1782; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1784 = 10'h29b == EXMEMALUOut[9:0] ? DMemory_667 : _GEN_1783; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1785 = 10'h29c == EXMEMALUOut[9:0] ? DMemory_668 : _GEN_1784; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1786 = 10'h29d == EXMEMALUOut[9:0] ? DMemory_669 : _GEN_1785; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1787 = 10'h29e == EXMEMALUOut[9:0] ? DMemory_670 : _GEN_1786; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1788 = 10'h29f == EXMEMALUOut[9:0] ? DMemory_671 : _GEN_1787; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1789 = 10'h2a0 == EXMEMALUOut[9:0] ? DMemory_672 : _GEN_1788; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1790 = 10'h2a1 == EXMEMALUOut[9:0] ? DMemory_673 : _GEN_1789; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1791 = 10'h2a2 == EXMEMALUOut[9:0] ? DMemory_674 : _GEN_1790; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1792 = 10'h2a3 == EXMEMALUOut[9:0] ? DMemory_675 : _GEN_1791; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1793 = 10'h2a4 == EXMEMALUOut[9:0] ? DMemory_676 : _GEN_1792; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1794 = 10'h2a5 == EXMEMALUOut[9:0] ? DMemory_677 : _GEN_1793; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1795 = 10'h2a6 == EXMEMALUOut[9:0] ? DMemory_678 : _GEN_1794; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1796 = 10'h2a7 == EXMEMALUOut[9:0] ? DMemory_679 : _GEN_1795; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1797 = 10'h2a8 == EXMEMALUOut[9:0] ? DMemory_680 : _GEN_1796; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1798 = 10'h2a9 == EXMEMALUOut[9:0] ? DMemory_681 : _GEN_1797; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1799 = 10'h2aa == EXMEMALUOut[9:0] ? DMemory_682 : _GEN_1798; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1800 = 10'h2ab == EXMEMALUOut[9:0] ? DMemory_683 : _GEN_1799; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1801 = 10'h2ac == EXMEMALUOut[9:0] ? DMemory_684 : _GEN_1800; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1802 = 10'h2ad == EXMEMALUOut[9:0] ? DMemory_685 : _GEN_1801; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1803 = 10'h2ae == EXMEMALUOut[9:0] ? DMemory_686 : _GEN_1802; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1804 = 10'h2af == EXMEMALUOut[9:0] ? DMemory_687 : _GEN_1803; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1805 = 10'h2b0 == EXMEMALUOut[9:0] ? DMemory_688 : _GEN_1804; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1806 = 10'h2b1 == EXMEMALUOut[9:0] ? DMemory_689 : _GEN_1805; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1807 = 10'h2b2 == EXMEMALUOut[9:0] ? DMemory_690 : _GEN_1806; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1808 = 10'h2b3 == EXMEMALUOut[9:0] ? DMemory_691 : _GEN_1807; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1809 = 10'h2b4 == EXMEMALUOut[9:0] ? DMemory_692 : _GEN_1808; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1810 = 10'h2b5 == EXMEMALUOut[9:0] ? DMemory_693 : _GEN_1809; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1811 = 10'h2b6 == EXMEMALUOut[9:0] ? DMemory_694 : _GEN_1810; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1812 = 10'h2b7 == EXMEMALUOut[9:0] ? DMemory_695 : _GEN_1811; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1813 = 10'h2b8 == EXMEMALUOut[9:0] ? DMemory_696 : _GEN_1812; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1814 = 10'h2b9 == EXMEMALUOut[9:0] ? DMemory_697 : _GEN_1813; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1815 = 10'h2ba == EXMEMALUOut[9:0] ? DMemory_698 : _GEN_1814; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1816 = 10'h2bb == EXMEMALUOut[9:0] ? DMemory_699 : _GEN_1815; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1817 = 10'h2bc == EXMEMALUOut[9:0] ? DMemory_700 : _GEN_1816; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1818 = 10'h2bd == EXMEMALUOut[9:0] ? DMemory_701 : _GEN_1817; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1819 = 10'h2be == EXMEMALUOut[9:0] ? DMemory_702 : _GEN_1818; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1820 = 10'h2bf == EXMEMALUOut[9:0] ? DMemory_703 : _GEN_1819; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1821 = 10'h2c0 == EXMEMALUOut[9:0] ? DMemory_704 : _GEN_1820; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1822 = 10'h2c1 == EXMEMALUOut[9:0] ? DMemory_705 : _GEN_1821; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1823 = 10'h2c2 == EXMEMALUOut[9:0] ? DMemory_706 : _GEN_1822; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1824 = 10'h2c3 == EXMEMALUOut[9:0] ? DMemory_707 : _GEN_1823; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1825 = 10'h2c4 == EXMEMALUOut[9:0] ? DMemory_708 : _GEN_1824; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1826 = 10'h2c5 == EXMEMALUOut[9:0] ? DMemory_709 : _GEN_1825; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1827 = 10'h2c6 == EXMEMALUOut[9:0] ? DMemory_710 : _GEN_1826; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1828 = 10'h2c7 == EXMEMALUOut[9:0] ? DMemory_711 : _GEN_1827; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1829 = 10'h2c8 == EXMEMALUOut[9:0] ? DMemory_712 : _GEN_1828; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1830 = 10'h2c9 == EXMEMALUOut[9:0] ? DMemory_713 : _GEN_1829; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1831 = 10'h2ca == EXMEMALUOut[9:0] ? DMemory_714 : _GEN_1830; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1832 = 10'h2cb == EXMEMALUOut[9:0] ? DMemory_715 : _GEN_1831; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1833 = 10'h2cc == EXMEMALUOut[9:0] ? DMemory_716 : _GEN_1832; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1834 = 10'h2cd == EXMEMALUOut[9:0] ? DMemory_717 : _GEN_1833; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1835 = 10'h2ce == EXMEMALUOut[9:0] ? DMemory_718 : _GEN_1834; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1836 = 10'h2cf == EXMEMALUOut[9:0] ? DMemory_719 : _GEN_1835; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1837 = 10'h2d0 == EXMEMALUOut[9:0] ? DMemory_720 : _GEN_1836; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1838 = 10'h2d1 == EXMEMALUOut[9:0] ? DMemory_721 : _GEN_1837; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1839 = 10'h2d2 == EXMEMALUOut[9:0] ? DMemory_722 : _GEN_1838; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1840 = 10'h2d3 == EXMEMALUOut[9:0] ? DMemory_723 : _GEN_1839; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1841 = 10'h2d4 == EXMEMALUOut[9:0] ? DMemory_724 : _GEN_1840; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1842 = 10'h2d5 == EXMEMALUOut[9:0] ? DMemory_725 : _GEN_1841; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1843 = 10'h2d6 == EXMEMALUOut[9:0] ? DMemory_726 : _GEN_1842; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1844 = 10'h2d7 == EXMEMALUOut[9:0] ? DMemory_727 : _GEN_1843; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1845 = 10'h2d8 == EXMEMALUOut[9:0] ? DMemory_728 : _GEN_1844; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1846 = 10'h2d9 == EXMEMALUOut[9:0] ? DMemory_729 : _GEN_1845; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1847 = 10'h2da == EXMEMALUOut[9:0] ? DMemory_730 : _GEN_1846; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1848 = 10'h2db == EXMEMALUOut[9:0] ? DMemory_731 : _GEN_1847; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1849 = 10'h2dc == EXMEMALUOut[9:0] ? DMemory_732 : _GEN_1848; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1850 = 10'h2dd == EXMEMALUOut[9:0] ? DMemory_733 : _GEN_1849; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1851 = 10'h2de == EXMEMALUOut[9:0] ? DMemory_734 : _GEN_1850; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1852 = 10'h2df == EXMEMALUOut[9:0] ? DMemory_735 : _GEN_1851; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1853 = 10'h2e0 == EXMEMALUOut[9:0] ? DMemory_736 : _GEN_1852; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1854 = 10'h2e1 == EXMEMALUOut[9:0] ? DMemory_737 : _GEN_1853; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1855 = 10'h2e2 == EXMEMALUOut[9:0] ? DMemory_738 : _GEN_1854; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1856 = 10'h2e3 == EXMEMALUOut[9:0] ? DMemory_739 : _GEN_1855; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1857 = 10'h2e4 == EXMEMALUOut[9:0] ? DMemory_740 : _GEN_1856; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1858 = 10'h2e5 == EXMEMALUOut[9:0] ? DMemory_741 : _GEN_1857; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1859 = 10'h2e6 == EXMEMALUOut[9:0] ? DMemory_742 : _GEN_1858; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1860 = 10'h2e7 == EXMEMALUOut[9:0] ? DMemory_743 : _GEN_1859; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1861 = 10'h2e8 == EXMEMALUOut[9:0] ? DMemory_744 : _GEN_1860; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1862 = 10'h2e9 == EXMEMALUOut[9:0] ? DMemory_745 : _GEN_1861; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1863 = 10'h2ea == EXMEMALUOut[9:0] ? DMemory_746 : _GEN_1862; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1864 = 10'h2eb == EXMEMALUOut[9:0] ? DMemory_747 : _GEN_1863; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1865 = 10'h2ec == EXMEMALUOut[9:0] ? DMemory_748 : _GEN_1864; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1866 = 10'h2ed == EXMEMALUOut[9:0] ? DMemory_749 : _GEN_1865; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1867 = 10'h2ee == EXMEMALUOut[9:0] ? DMemory_750 : _GEN_1866; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1868 = 10'h2ef == EXMEMALUOut[9:0] ? DMemory_751 : _GEN_1867; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1869 = 10'h2f0 == EXMEMALUOut[9:0] ? DMemory_752 : _GEN_1868; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1870 = 10'h2f1 == EXMEMALUOut[9:0] ? DMemory_753 : _GEN_1869; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1871 = 10'h2f2 == EXMEMALUOut[9:0] ? DMemory_754 : _GEN_1870; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1872 = 10'h2f3 == EXMEMALUOut[9:0] ? DMemory_755 : _GEN_1871; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1873 = 10'h2f4 == EXMEMALUOut[9:0] ? DMemory_756 : _GEN_1872; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1874 = 10'h2f5 == EXMEMALUOut[9:0] ? DMemory_757 : _GEN_1873; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1875 = 10'h2f6 == EXMEMALUOut[9:0] ? DMemory_758 : _GEN_1874; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1876 = 10'h2f7 == EXMEMALUOut[9:0] ? DMemory_759 : _GEN_1875; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1877 = 10'h2f8 == EXMEMALUOut[9:0] ? DMemory_760 : _GEN_1876; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1878 = 10'h2f9 == EXMEMALUOut[9:0] ? DMemory_761 : _GEN_1877; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1879 = 10'h2fa == EXMEMALUOut[9:0] ? DMemory_762 : _GEN_1878; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1880 = 10'h2fb == EXMEMALUOut[9:0] ? DMemory_763 : _GEN_1879; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1881 = 10'h2fc == EXMEMALUOut[9:0] ? DMemory_764 : _GEN_1880; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1882 = 10'h2fd == EXMEMALUOut[9:0] ? DMemory_765 : _GEN_1881; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1883 = 10'h2fe == EXMEMALUOut[9:0] ? DMemory_766 : _GEN_1882; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1884 = 10'h2ff == EXMEMALUOut[9:0] ? DMemory_767 : _GEN_1883; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1885 = 10'h300 == EXMEMALUOut[9:0] ? DMemory_768 : _GEN_1884; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1886 = 10'h301 == EXMEMALUOut[9:0] ? DMemory_769 : _GEN_1885; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1887 = 10'h302 == EXMEMALUOut[9:0] ? DMemory_770 : _GEN_1886; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1888 = 10'h303 == EXMEMALUOut[9:0] ? DMemory_771 : _GEN_1887; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1889 = 10'h304 == EXMEMALUOut[9:0] ? DMemory_772 : _GEN_1888; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1890 = 10'h305 == EXMEMALUOut[9:0] ? DMemory_773 : _GEN_1889; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1891 = 10'h306 == EXMEMALUOut[9:0] ? DMemory_774 : _GEN_1890; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1892 = 10'h307 == EXMEMALUOut[9:0] ? DMemory_775 : _GEN_1891; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1893 = 10'h308 == EXMEMALUOut[9:0] ? DMemory_776 : _GEN_1892; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1894 = 10'h309 == EXMEMALUOut[9:0] ? DMemory_777 : _GEN_1893; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1895 = 10'h30a == EXMEMALUOut[9:0] ? DMemory_778 : _GEN_1894; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1896 = 10'h30b == EXMEMALUOut[9:0] ? DMemory_779 : _GEN_1895; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1897 = 10'h30c == EXMEMALUOut[9:0] ? DMemory_780 : _GEN_1896; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1898 = 10'h30d == EXMEMALUOut[9:0] ? DMemory_781 : _GEN_1897; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1899 = 10'h30e == EXMEMALUOut[9:0] ? DMemory_782 : _GEN_1898; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1900 = 10'h30f == EXMEMALUOut[9:0] ? DMemory_783 : _GEN_1899; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1901 = 10'h310 == EXMEMALUOut[9:0] ? DMemory_784 : _GEN_1900; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1902 = 10'h311 == EXMEMALUOut[9:0] ? DMemory_785 : _GEN_1901; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1903 = 10'h312 == EXMEMALUOut[9:0] ? DMemory_786 : _GEN_1902; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1904 = 10'h313 == EXMEMALUOut[9:0] ? DMemory_787 : _GEN_1903; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1905 = 10'h314 == EXMEMALUOut[9:0] ? DMemory_788 : _GEN_1904; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1906 = 10'h315 == EXMEMALUOut[9:0] ? DMemory_789 : _GEN_1905; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1907 = 10'h316 == EXMEMALUOut[9:0] ? DMemory_790 : _GEN_1906; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1908 = 10'h317 == EXMEMALUOut[9:0] ? DMemory_791 : _GEN_1907; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1909 = 10'h318 == EXMEMALUOut[9:0] ? DMemory_792 : _GEN_1908; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1910 = 10'h319 == EXMEMALUOut[9:0] ? DMemory_793 : _GEN_1909; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1911 = 10'h31a == EXMEMALUOut[9:0] ? DMemory_794 : _GEN_1910; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1912 = 10'h31b == EXMEMALUOut[9:0] ? DMemory_795 : _GEN_1911; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1913 = 10'h31c == EXMEMALUOut[9:0] ? DMemory_796 : _GEN_1912; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1914 = 10'h31d == EXMEMALUOut[9:0] ? DMemory_797 : _GEN_1913; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1915 = 10'h31e == EXMEMALUOut[9:0] ? DMemory_798 : _GEN_1914; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1916 = 10'h31f == EXMEMALUOut[9:0] ? DMemory_799 : _GEN_1915; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1917 = 10'h320 == EXMEMALUOut[9:0] ? DMemory_800 : _GEN_1916; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1918 = 10'h321 == EXMEMALUOut[9:0] ? DMemory_801 : _GEN_1917; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1919 = 10'h322 == EXMEMALUOut[9:0] ? DMemory_802 : _GEN_1918; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1920 = 10'h323 == EXMEMALUOut[9:0] ? DMemory_803 : _GEN_1919; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1921 = 10'h324 == EXMEMALUOut[9:0] ? DMemory_804 : _GEN_1920; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1922 = 10'h325 == EXMEMALUOut[9:0] ? DMemory_805 : _GEN_1921; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1923 = 10'h326 == EXMEMALUOut[9:0] ? DMemory_806 : _GEN_1922; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1924 = 10'h327 == EXMEMALUOut[9:0] ? DMemory_807 : _GEN_1923; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1925 = 10'h328 == EXMEMALUOut[9:0] ? DMemory_808 : _GEN_1924; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1926 = 10'h329 == EXMEMALUOut[9:0] ? DMemory_809 : _GEN_1925; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1927 = 10'h32a == EXMEMALUOut[9:0] ? DMemory_810 : _GEN_1926; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1928 = 10'h32b == EXMEMALUOut[9:0] ? DMemory_811 : _GEN_1927; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1929 = 10'h32c == EXMEMALUOut[9:0] ? DMemory_812 : _GEN_1928; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1930 = 10'h32d == EXMEMALUOut[9:0] ? DMemory_813 : _GEN_1929; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1931 = 10'h32e == EXMEMALUOut[9:0] ? DMemory_814 : _GEN_1930; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1932 = 10'h32f == EXMEMALUOut[9:0] ? DMemory_815 : _GEN_1931; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1933 = 10'h330 == EXMEMALUOut[9:0] ? DMemory_816 : _GEN_1932; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1934 = 10'h331 == EXMEMALUOut[9:0] ? DMemory_817 : _GEN_1933; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1935 = 10'h332 == EXMEMALUOut[9:0] ? DMemory_818 : _GEN_1934; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1936 = 10'h333 == EXMEMALUOut[9:0] ? DMemory_819 : _GEN_1935; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1937 = 10'h334 == EXMEMALUOut[9:0] ? DMemory_820 : _GEN_1936; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1938 = 10'h335 == EXMEMALUOut[9:0] ? DMemory_821 : _GEN_1937; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1939 = 10'h336 == EXMEMALUOut[9:0] ? DMemory_822 : _GEN_1938; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1940 = 10'h337 == EXMEMALUOut[9:0] ? DMemory_823 : _GEN_1939; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1941 = 10'h338 == EXMEMALUOut[9:0] ? DMemory_824 : _GEN_1940; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1942 = 10'h339 == EXMEMALUOut[9:0] ? DMemory_825 : _GEN_1941; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1943 = 10'h33a == EXMEMALUOut[9:0] ? DMemory_826 : _GEN_1942; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1944 = 10'h33b == EXMEMALUOut[9:0] ? DMemory_827 : _GEN_1943; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1945 = 10'h33c == EXMEMALUOut[9:0] ? DMemory_828 : _GEN_1944; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1946 = 10'h33d == EXMEMALUOut[9:0] ? DMemory_829 : _GEN_1945; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1947 = 10'h33e == EXMEMALUOut[9:0] ? DMemory_830 : _GEN_1946; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1948 = 10'h33f == EXMEMALUOut[9:0] ? DMemory_831 : _GEN_1947; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1949 = 10'h340 == EXMEMALUOut[9:0] ? DMemory_832 : _GEN_1948; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1950 = 10'h341 == EXMEMALUOut[9:0] ? DMemory_833 : _GEN_1949; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1951 = 10'h342 == EXMEMALUOut[9:0] ? DMemory_834 : _GEN_1950; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1952 = 10'h343 == EXMEMALUOut[9:0] ? DMemory_835 : _GEN_1951; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1953 = 10'h344 == EXMEMALUOut[9:0] ? DMemory_836 : _GEN_1952; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1954 = 10'h345 == EXMEMALUOut[9:0] ? DMemory_837 : _GEN_1953; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1955 = 10'h346 == EXMEMALUOut[9:0] ? DMemory_838 : _GEN_1954; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1956 = 10'h347 == EXMEMALUOut[9:0] ? DMemory_839 : _GEN_1955; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1957 = 10'h348 == EXMEMALUOut[9:0] ? DMemory_840 : _GEN_1956; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1958 = 10'h349 == EXMEMALUOut[9:0] ? DMemory_841 : _GEN_1957; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1959 = 10'h34a == EXMEMALUOut[9:0] ? DMemory_842 : _GEN_1958; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1960 = 10'h34b == EXMEMALUOut[9:0] ? DMemory_843 : _GEN_1959; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1961 = 10'h34c == EXMEMALUOut[9:0] ? DMemory_844 : _GEN_1960; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1962 = 10'h34d == EXMEMALUOut[9:0] ? DMemory_845 : _GEN_1961; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1963 = 10'h34e == EXMEMALUOut[9:0] ? DMemory_846 : _GEN_1962; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1964 = 10'h34f == EXMEMALUOut[9:0] ? DMemory_847 : _GEN_1963; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1965 = 10'h350 == EXMEMALUOut[9:0] ? DMemory_848 : _GEN_1964; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1966 = 10'h351 == EXMEMALUOut[9:0] ? DMemory_849 : _GEN_1965; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1967 = 10'h352 == EXMEMALUOut[9:0] ? DMemory_850 : _GEN_1966; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1968 = 10'h353 == EXMEMALUOut[9:0] ? DMemory_851 : _GEN_1967; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1969 = 10'h354 == EXMEMALUOut[9:0] ? DMemory_852 : _GEN_1968; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1970 = 10'h355 == EXMEMALUOut[9:0] ? DMemory_853 : _GEN_1969; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1971 = 10'h356 == EXMEMALUOut[9:0] ? DMemory_854 : _GEN_1970; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1972 = 10'h357 == EXMEMALUOut[9:0] ? DMemory_855 : _GEN_1971; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1973 = 10'h358 == EXMEMALUOut[9:0] ? DMemory_856 : _GEN_1972; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1974 = 10'h359 == EXMEMALUOut[9:0] ? DMemory_857 : _GEN_1973; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1975 = 10'h35a == EXMEMALUOut[9:0] ? DMemory_858 : _GEN_1974; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1976 = 10'h35b == EXMEMALUOut[9:0] ? DMemory_859 : _GEN_1975; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1977 = 10'h35c == EXMEMALUOut[9:0] ? DMemory_860 : _GEN_1976; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1978 = 10'h35d == EXMEMALUOut[9:0] ? DMemory_861 : _GEN_1977; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1979 = 10'h35e == EXMEMALUOut[9:0] ? DMemory_862 : _GEN_1978; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1980 = 10'h35f == EXMEMALUOut[9:0] ? DMemory_863 : _GEN_1979; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1981 = 10'h360 == EXMEMALUOut[9:0] ? DMemory_864 : _GEN_1980; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1982 = 10'h361 == EXMEMALUOut[9:0] ? DMemory_865 : _GEN_1981; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1983 = 10'h362 == EXMEMALUOut[9:0] ? DMemory_866 : _GEN_1982; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1984 = 10'h363 == EXMEMALUOut[9:0] ? DMemory_867 : _GEN_1983; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1985 = 10'h364 == EXMEMALUOut[9:0] ? DMemory_868 : _GEN_1984; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1986 = 10'h365 == EXMEMALUOut[9:0] ? DMemory_869 : _GEN_1985; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1987 = 10'h366 == EXMEMALUOut[9:0] ? DMemory_870 : _GEN_1986; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1988 = 10'h367 == EXMEMALUOut[9:0] ? DMemory_871 : _GEN_1987; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1989 = 10'h368 == EXMEMALUOut[9:0] ? DMemory_872 : _GEN_1988; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1990 = 10'h369 == EXMEMALUOut[9:0] ? DMemory_873 : _GEN_1989; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1991 = 10'h36a == EXMEMALUOut[9:0] ? DMemory_874 : _GEN_1990; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1992 = 10'h36b == EXMEMALUOut[9:0] ? DMemory_875 : _GEN_1991; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1993 = 10'h36c == EXMEMALUOut[9:0] ? DMemory_876 : _GEN_1992; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1994 = 10'h36d == EXMEMALUOut[9:0] ? DMemory_877 : _GEN_1993; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1995 = 10'h36e == EXMEMALUOut[9:0] ? DMemory_878 : _GEN_1994; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1996 = 10'h36f == EXMEMALUOut[9:0] ? DMemory_879 : _GEN_1995; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1997 = 10'h370 == EXMEMALUOut[9:0] ? DMemory_880 : _GEN_1996; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1998 = 10'h371 == EXMEMALUOut[9:0] ? DMemory_881 : _GEN_1997; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_1999 = 10'h372 == EXMEMALUOut[9:0] ? DMemory_882 : _GEN_1998; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2000 = 10'h373 == EXMEMALUOut[9:0] ? DMemory_883 : _GEN_1999; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2001 = 10'h374 == EXMEMALUOut[9:0] ? DMemory_884 : _GEN_2000; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2002 = 10'h375 == EXMEMALUOut[9:0] ? DMemory_885 : _GEN_2001; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2003 = 10'h376 == EXMEMALUOut[9:0] ? DMemory_886 : _GEN_2002; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2004 = 10'h377 == EXMEMALUOut[9:0] ? DMemory_887 : _GEN_2003; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2005 = 10'h378 == EXMEMALUOut[9:0] ? DMemory_888 : _GEN_2004; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2006 = 10'h379 == EXMEMALUOut[9:0] ? DMemory_889 : _GEN_2005; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2007 = 10'h37a == EXMEMALUOut[9:0] ? DMemory_890 : _GEN_2006; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2008 = 10'h37b == EXMEMALUOut[9:0] ? DMemory_891 : _GEN_2007; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2009 = 10'h37c == EXMEMALUOut[9:0] ? DMemory_892 : _GEN_2008; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2010 = 10'h37d == EXMEMALUOut[9:0] ? DMemory_893 : _GEN_2009; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2011 = 10'h37e == EXMEMALUOut[9:0] ? DMemory_894 : _GEN_2010; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2012 = 10'h37f == EXMEMALUOut[9:0] ? DMemory_895 : _GEN_2011; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2013 = 10'h380 == EXMEMALUOut[9:0] ? DMemory_896 : _GEN_2012; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2014 = 10'h381 == EXMEMALUOut[9:0] ? DMemory_897 : _GEN_2013; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2015 = 10'h382 == EXMEMALUOut[9:0] ? DMemory_898 : _GEN_2014; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2016 = 10'h383 == EXMEMALUOut[9:0] ? DMemory_899 : _GEN_2015; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2017 = 10'h384 == EXMEMALUOut[9:0] ? DMemory_900 : _GEN_2016; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2018 = 10'h385 == EXMEMALUOut[9:0] ? DMemory_901 : _GEN_2017; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2019 = 10'h386 == EXMEMALUOut[9:0] ? DMemory_902 : _GEN_2018; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2020 = 10'h387 == EXMEMALUOut[9:0] ? DMemory_903 : _GEN_2019; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2021 = 10'h388 == EXMEMALUOut[9:0] ? DMemory_904 : _GEN_2020; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2022 = 10'h389 == EXMEMALUOut[9:0] ? DMemory_905 : _GEN_2021; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2023 = 10'h38a == EXMEMALUOut[9:0] ? DMemory_906 : _GEN_2022; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2024 = 10'h38b == EXMEMALUOut[9:0] ? DMemory_907 : _GEN_2023; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2025 = 10'h38c == EXMEMALUOut[9:0] ? DMemory_908 : _GEN_2024; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2026 = 10'h38d == EXMEMALUOut[9:0] ? DMemory_909 : _GEN_2025; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2027 = 10'h38e == EXMEMALUOut[9:0] ? DMemory_910 : _GEN_2026; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2028 = 10'h38f == EXMEMALUOut[9:0] ? DMemory_911 : _GEN_2027; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2029 = 10'h390 == EXMEMALUOut[9:0] ? DMemory_912 : _GEN_2028; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2030 = 10'h391 == EXMEMALUOut[9:0] ? DMemory_913 : _GEN_2029; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2031 = 10'h392 == EXMEMALUOut[9:0] ? DMemory_914 : _GEN_2030; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2032 = 10'h393 == EXMEMALUOut[9:0] ? DMemory_915 : _GEN_2031; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2033 = 10'h394 == EXMEMALUOut[9:0] ? DMemory_916 : _GEN_2032; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2034 = 10'h395 == EXMEMALUOut[9:0] ? DMemory_917 : _GEN_2033; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2035 = 10'h396 == EXMEMALUOut[9:0] ? DMemory_918 : _GEN_2034; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2036 = 10'h397 == EXMEMALUOut[9:0] ? DMemory_919 : _GEN_2035; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2037 = 10'h398 == EXMEMALUOut[9:0] ? DMemory_920 : _GEN_2036; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2038 = 10'h399 == EXMEMALUOut[9:0] ? DMemory_921 : _GEN_2037; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2039 = 10'h39a == EXMEMALUOut[9:0] ? DMemory_922 : _GEN_2038; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2040 = 10'h39b == EXMEMALUOut[9:0] ? DMemory_923 : _GEN_2039; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2041 = 10'h39c == EXMEMALUOut[9:0] ? DMemory_924 : _GEN_2040; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2042 = 10'h39d == EXMEMALUOut[9:0] ? DMemory_925 : _GEN_2041; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2043 = 10'h39e == EXMEMALUOut[9:0] ? DMemory_926 : _GEN_2042; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2044 = 10'h39f == EXMEMALUOut[9:0] ? DMemory_927 : _GEN_2043; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2045 = 10'h3a0 == EXMEMALUOut[9:0] ? DMemory_928 : _GEN_2044; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2046 = 10'h3a1 == EXMEMALUOut[9:0] ? DMemory_929 : _GEN_2045; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2047 = 10'h3a2 == EXMEMALUOut[9:0] ? DMemory_930 : _GEN_2046; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2048 = 10'h3a3 == EXMEMALUOut[9:0] ? DMemory_931 : _GEN_2047; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2049 = 10'h3a4 == EXMEMALUOut[9:0] ? DMemory_932 : _GEN_2048; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2050 = 10'h3a5 == EXMEMALUOut[9:0] ? DMemory_933 : _GEN_2049; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2051 = 10'h3a6 == EXMEMALUOut[9:0] ? DMemory_934 : _GEN_2050; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2052 = 10'h3a7 == EXMEMALUOut[9:0] ? DMemory_935 : _GEN_2051; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2053 = 10'h3a8 == EXMEMALUOut[9:0] ? DMemory_936 : _GEN_2052; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2054 = 10'h3a9 == EXMEMALUOut[9:0] ? DMemory_937 : _GEN_2053; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2055 = 10'h3aa == EXMEMALUOut[9:0] ? DMemory_938 : _GEN_2054; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2056 = 10'h3ab == EXMEMALUOut[9:0] ? DMemory_939 : _GEN_2055; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2057 = 10'h3ac == EXMEMALUOut[9:0] ? DMemory_940 : _GEN_2056; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2058 = 10'h3ad == EXMEMALUOut[9:0] ? DMemory_941 : _GEN_2057; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2059 = 10'h3ae == EXMEMALUOut[9:0] ? DMemory_942 : _GEN_2058; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2060 = 10'h3af == EXMEMALUOut[9:0] ? DMemory_943 : _GEN_2059; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2061 = 10'h3b0 == EXMEMALUOut[9:0] ? DMemory_944 : _GEN_2060; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2062 = 10'h3b1 == EXMEMALUOut[9:0] ? DMemory_945 : _GEN_2061; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2063 = 10'h3b2 == EXMEMALUOut[9:0] ? DMemory_946 : _GEN_2062; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2064 = 10'h3b3 == EXMEMALUOut[9:0] ? DMemory_947 : _GEN_2063; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2065 = 10'h3b4 == EXMEMALUOut[9:0] ? DMemory_948 : _GEN_2064; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2066 = 10'h3b5 == EXMEMALUOut[9:0] ? DMemory_949 : _GEN_2065; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2067 = 10'h3b6 == EXMEMALUOut[9:0] ? DMemory_950 : _GEN_2066; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2068 = 10'h3b7 == EXMEMALUOut[9:0] ? DMemory_951 : _GEN_2067; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2069 = 10'h3b8 == EXMEMALUOut[9:0] ? DMemory_952 : _GEN_2068; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2070 = 10'h3b9 == EXMEMALUOut[9:0] ? DMemory_953 : _GEN_2069; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2071 = 10'h3ba == EXMEMALUOut[9:0] ? DMemory_954 : _GEN_2070; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2072 = 10'h3bb == EXMEMALUOut[9:0] ? DMemory_955 : _GEN_2071; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2073 = 10'h3bc == EXMEMALUOut[9:0] ? DMemory_956 : _GEN_2072; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2074 = 10'h3bd == EXMEMALUOut[9:0] ? DMemory_957 : _GEN_2073; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2075 = 10'h3be == EXMEMALUOut[9:0] ? DMemory_958 : _GEN_2074; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2076 = 10'h3bf == EXMEMALUOut[9:0] ? DMemory_959 : _GEN_2075; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2077 = 10'h3c0 == EXMEMALUOut[9:0] ? DMemory_960 : _GEN_2076; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2078 = 10'h3c1 == EXMEMALUOut[9:0] ? DMemory_961 : _GEN_2077; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2079 = 10'h3c2 == EXMEMALUOut[9:0] ? DMemory_962 : _GEN_2078; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2080 = 10'h3c3 == EXMEMALUOut[9:0] ? DMemory_963 : _GEN_2079; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2081 = 10'h3c4 == EXMEMALUOut[9:0] ? DMemory_964 : _GEN_2080; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2082 = 10'h3c5 == EXMEMALUOut[9:0] ? DMemory_965 : _GEN_2081; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2083 = 10'h3c6 == EXMEMALUOut[9:0] ? DMemory_966 : _GEN_2082; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2084 = 10'h3c7 == EXMEMALUOut[9:0] ? DMemory_967 : _GEN_2083; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2085 = 10'h3c8 == EXMEMALUOut[9:0] ? DMemory_968 : _GEN_2084; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2086 = 10'h3c9 == EXMEMALUOut[9:0] ? DMemory_969 : _GEN_2085; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2087 = 10'h3ca == EXMEMALUOut[9:0] ? DMemory_970 : _GEN_2086; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2088 = 10'h3cb == EXMEMALUOut[9:0] ? DMemory_971 : _GEN_2087; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2089 = 10'h3cc == EXMEMALUOut[9:0] ? DMemory_972 : _GEN_2088; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2090 = 10'h3cd == EXMEMALUOut[9:0] ? DMemory_973 : _GEN_2089; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2091 = 10'h3ce == EXMEMALUOut[9:0] ? DMemory_974 : _GEN_2090; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2092 = 10'h3cf == EXMEMALUOut[9:0] ? DMemory_975 : _GEN_2091; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2093 = 10'h3d0 == EXMEMALUOut[9:0] ? DMemory_976 : _GEN_2092; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2094 = 10'h3d1 == EXMEMALUOut[9:0] ? DMemory_977 : _GEN_2093; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2095 = 10'h3d2 == EXMEMALUOut[9:0] ? DMemory_978 : _GEN_2094; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2096 = 10'h3d3 == EXMEMALUOut[9:0] ? DMemory_979 : _GEN_2095; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2097 = 10'h3d4 == EXMEMALUOut[9:0] ? DMemory_980 : _GEN_2096; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2098 = 10'h3d5 == EXMEMALUOut[9:0] ? DMemory_981 : _GEN_2097; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2099 = 10'h3d6 == EXMEMALUOut[9:0] ? DMemory_982 : _GEN_2098; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2100 = 10'h3d7 == EXMEMALUOut[9:0] ? DMemory_983 : _GEN_2099; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2101 = 10'h3d8 == EXMEMALUOut[9:0] ? DMemory_984 : _GEN_2100; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2102 = 10'h3d9 == EXMEMALUOut[9:0] ? DMemory_985 : _GEN_2101; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2103 = 10'h3da == EXMEMALUOut[9:0] ? DMemory_986 : _GEN_2102; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2104 = 10'h3db == EXMEMALUOut[9:0] ? DMemory_987 : _GEN_2103; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2105 = 10'h3dc == EXMEMALUOut[9:0] ? DMemory_988 : _GEN_2104; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2106 = 10'h3dd == EXMEMALUOut[9:0] ? DMemory_989 : _GEN_2105; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2107 = 10'h3de == EXMEMALUOut[9:0] ? DMemory_990 : _GEN_2106; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2108 = 10'h3df == EXMEMALUOut[9:0] ? DMemory_991 : _GEN_2107; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2109 = 10'h3e0 == EXMEMALUOut[9:0] ? DMemory_992 : _GEN_2108; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2110 = 10'h3e1 == EXMEMALUOut[9:0] ? DMemory_993 : _GEN_2109; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2111 = 10'h3e2 == EXMEMALUOut[9:0] ? DMemory_994 : _GEN_2110; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2112 = 10'h3e3 == EXMEMALUOut[9:0] ? DMemory_995 : _GEN_2111; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2113 = 10'h3e4 == EXMEMALUOut[9:0] ? DMemory_996 : _GEN_2112; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2114 = 10'h3e5 == EXMEMALUOut[9:0] ? DMemory_997 : _GEN_2113; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2115 = 10'h3e6 == EXMEMALUOut[9:0] ? DMemory_998 : _GEN_2114; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2116 = 10'h3e7 == EXMEMALUOut[9:0] ? DMemory_999 : _GEN_2115; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2117 = 10'h3e8 == EXMEMALUOut[9:0] ? DMemory_1000 : _GEN_2116; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2118 = 10'h3e9 == EXMEMALUOut[9:0] ? DMemory_1001 : _GEN_2117; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2119 = 10'h3ea == EXMEMALUOut[9:0] ? DMemory_1002 : _GEN_2118; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2120 = 10'h3eb == EXMEMALUOut[9:0] ? DMemory_1003 : _GEN_2119; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2121 = 10'h3ec == EXMEMALUOut[9:0] ? DMemory_1004 : _GEN_2120; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2122 = 10'h3ed == EXMEMALUOut[9:0] ? DMemory_1005 : _GEN_2121; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2123 = 10'h3ee == EXMEMALUOut[9:0] ? DMemory_1006 : _GEN_2122; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2124 = 10'h3ef == EXMEMALUOut[9:0] ? DMemory_1007 : _GEN_2123; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2125 = 10'h3f0 == EXMEMALUOut[9:0] ? DMemory_1008 : _GEN_2124; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2126 = 10'h3f1 == EXMEMALUOut[9:0] ? DMemory_1009 : _GEN_2125; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2127 = 10'h3f2 == EXMEMALUOut[9:0] ? DMemory_1010 : _GEN_2126; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2128 = 10'h3f3 == EXMEMALUOut[9:0] ? DMemory_1011 : _GEN_2127; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2129 = 10'h3f4 == EXMEMALUOut[9:0] ? DMemory_1012 : _GEN_2128; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2130 = 10'h3f5 == EXMEMALUOut[9:0] ? DMemory_1013 : _GEN_2129; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2131 = 10'h3f6 == EXMEMALUOut[9:0] ? DMemory_1014 : _GEN_2130; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2132 = 10'h3f7 == EXMEMALUOut[9:0] ? DMemory_1015 : _GEN_2131; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2133 = 10'h3f8 == EXMEMALUOut[9:0] ? DMemory_1016 : _GEN_2132; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2134 = 10'h3f9 == EXMEMALUOut[9:0] ? DMemory_1017 : _GEN_2133; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2135 = 10'h3fa == EXMEMALUOut[9:0] ? DMemory_1018 : _GEN_2134; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2136 = 10'h3fb == EXMEMALUOut[9:0] ? DMemory_1019 : _GEN_2135; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2137 = 10'h3fc == EXMEMALUOut[9:0] ? DMemory_1020 : _GEN_2136; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2138 = 10'h3fd == EXMEMALUOut[9:0] ? DMemory_1021 : _GEN_2137; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2139 = 10'h3fe == EXMEMALUOut[9:0] ? DMemory_1022 : _GEN_2138; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2140 = 10'h3ff == EXMEMALUOut[9:0] ? DMemory_1023 : _GEN_2139; // @[cpu.scala 219:{18,18}]
  wire [31:0] _GEN_2141 = 10'h0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_0; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2142 = 10'h1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2143 = 10'h2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_2; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2144 = 10'h3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_3; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2145 = 10'h4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_4; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2146 = 10'h5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_5; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2147 = 10'h6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_6; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2148 = 10'h7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_7; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2149 = 10'h8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_8; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2150 = 10'h9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_9; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2151 = 10'ha == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_10; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2152 = 10'hb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_11; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2153 = 10'hc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_12; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2154 = 10'hd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_13; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2155 = 10'he == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_14; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2156 = 10'hf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_15; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2157 = 10'h10 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_16; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2158 = 10'h11 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_17; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2159 = 10'h12 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_18; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2160 = 10'h13 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_19; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2161 = 10'h14 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_20; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2162 = 10'h15 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_21; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2163 = 10'h16 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_22; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2164 = 10'h17 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_23; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2165 = 10'h18 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_24; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2166 = 10'h19 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_25; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2167 = 10'h1a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_26; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2168 = 10'h1b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_27; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2169 = 10'h1c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_28; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2170 = 10'h1d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_29; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2171 = 10'h1e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_30; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2172 = 10'h1f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_31; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2173 = 10'h20 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_32; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2174 = 10'h21 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_33; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2175 = 10'h22 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_34; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2176 = 10'h23 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_35; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2177 = 10'h24 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_36; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2178 = 10'h25 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_37; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2179 = 10'h26 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_38; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2180 = 10'h27 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_39; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2181 = 10'h28 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_40; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2182 = 10'h29 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_41; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2183 = 10'h2a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_42; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2184 = 10'h2b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_43; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2185 = 10'h2c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_44; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2186 = 10'h2d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_45; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2187 = 10'h2e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_46; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2188 = 10'h2f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_47; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2189 = 10'h30 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_48; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2190 = 10'h31 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_49; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2191 = 10'h32 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_50; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2192 = 10'h33 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_51; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2193 = 10'h34 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_52; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2194 = 10'h35 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_53; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2195 = 10'h36 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_54; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2196 = 10'h37 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_55; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2197 = 10'h38 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_56; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2198 = 10'h39 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_57; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2199 = 10'h3a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_58; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2200 = 10'h3b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_59; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2201 = 10'h3c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_60; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2202 = 10'h3d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_61; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2203 = 10'h3e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_62; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2204 = 10'h3f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_63; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2205 = 10'h40 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_64; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2206 = 10'h41 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_65; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2207 = 10'h42 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_66; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2208 = 10'h43 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_67; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2209 = 10'h44 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_68; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2210 = 10'h45 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_69; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2211 = 10'h46 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_70; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2212 = 10'h47 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_71; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2213 = 10'h48 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_72; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2214 = 10'h49 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_73; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2215 = 10'h4a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_74; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2216 = 10'h4b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_75; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2217 = 10'h4c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_76; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2218 = 10'h4d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_77; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2219 = 10'h4e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_78; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2220 = 10'h4f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_79; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2221 = 10'h50 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_80; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2222 = 10'h51 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_81; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2223 = 10'h52 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_82; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2224 = 10'h53 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_83; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2225 = 10'h54 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_84; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2226 = 10'h55 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_85; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2227 = 10'h56 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_86; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2228 = 10'h57 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_87; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2229 = 10'h58 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_88; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2230 = 10'h59 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_89; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2231 = 10'h5a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_90; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2232 = 10'h5b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_91; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2233 = 10'h5c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_92; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2234 = 10'h5d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_93; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2235 = 10'h5e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_94; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2236 = 10'h5f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_95; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2237 = 10'h60 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_96; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2238 = 10'h61 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_97; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2239 = 10'h62 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_98; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2240 = 10'h63 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_99; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2241 = 10'h64 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_100; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2242 = 10'h65 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_101; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2243 = 10'h66 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_102; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2244 = 10'h67 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_103; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2245 = 10'h68 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_104; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2246 = 10'h69 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_105; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2247 = 10'h6a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_106; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2248 = 10'h6b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_107; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2249 = 10'h6c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_108; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2250 = 10'h6d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_109; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2251 = 10'h6e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_110; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2252 = 10'h6f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_111; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2253 = 10'h70 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_112; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2254 = 10'h71 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_113; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2255 = 10'h72 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_114; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2256 = 10'h73 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_115; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2257 = 10'h74 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_116; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2258 = 10'h75 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_117; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2259 = 10'h76 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_118; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2260 = 10'h77 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_119; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2261 = 10'h78 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_120; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2262 = 10'h79 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_121; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2263 = 10'h7a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_122; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2264 = 10'h7b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_123; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2265 = 10'h7c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_124; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2266 = 10'h7d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_125; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2267 = 10'h7e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_126; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2268 = 10'h7f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_127; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2269 = 10'h80 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_128; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2270 = 10'h81 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_129; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2271 = 10'h82 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_130; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2272 = 10'h83 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_131; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2273 = 10'h84 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_132; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2274 = 10'h85 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_133; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2275 = 10'h86 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_134; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2276 = 10'h87 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_135; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2277 = 10'h88 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_136; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2278 = 10'h89 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_137; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2279 = 10'h8a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_138; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2280 = 10'h8b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_139; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2281 = 10'h8c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_140; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2282 = 10'h8d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_141; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2283 = 10'h8e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_142; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2284 = 10'h8f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_143; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2285 = 10'h90 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_144; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2286 = 10'h91 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_145; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2287 = 10'h92 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_146; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2288 = 10'h93 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_147; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2289 = 10'h94 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_148; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2290 = 10'h95 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_149; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2291 = 10'h96 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_150; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2292 = 10'h97 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_151; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2293 = 10'h98 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_152; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2294 = 10'h99 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_153; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2295 = 10'h9a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_154; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2296 = 10'h9b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_155; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2297 = 10'h9c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_156; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2298 = 10'h9d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_157; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2299 = 10'h9e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_158; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2300 = 10'h9f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_159; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2301 = 10'ha0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_160; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2302 = 10'ha1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_161; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2303 = 10'ha2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_162; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2304 = 10'ha3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_163; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2305 = 10'ha4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_164; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2306 = 10'ha5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_165; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2307 = 10'ha6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_166; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2308 = 10'ha7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_167; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2309 = 10'ha8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_168; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2310 = 10'ha9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_169; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2311 = 10'haa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_170; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2312 = 10'hab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_171; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2313 = 10'hac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_172; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2314 = 10'had == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_173; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2315 = 10'hae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_174; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2316 = 10'haf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_175; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2317 = 10'hb0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_176; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2318 = 10'hb1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_177; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2319 = 10'hb2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_178; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2320 = 10'hb3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_179; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2321 = 10'hb4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_180; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2322 = 10'hb5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_181; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2323 = 10'hb6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_182; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2324 = 10'hb7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_183; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2325 = 10'hb8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_184; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2326 = 10'hb9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_185; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2327 = 10'hba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_186; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2328 = 10'hbb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_187; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2329 = 10'hbc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_188; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2330 = 10'hbd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_189; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2331 = 10'hbe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_190; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2332 = 10'hbf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_191; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2333 = 10'hc0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_192; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2334 = 10'hc1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_193; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2335 = 10'hc2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_194; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2336 = 10'hc3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_195; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2337 = 10'hc4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_196; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2338 = 10'hc5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_197; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2339 = 10'hc6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_198; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2340 = 10'hc7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_199; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2341 = 10'hc8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_200; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2342 = 10'hc9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_201; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2343 = 10'hca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_202; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2344 = 10'hcb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_203; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2345 = 10'hcc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_204; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2346 = 10'hcd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_205; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2347 = 10'hce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_206; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2348 = 10'hcf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_207; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2349 = 10'hd0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_208; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2350 = 10'hd1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_209; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2351 = 10'hd2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_210; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2352 = 10'hd3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_211; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2353 = 10'hd4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_212; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2354 = 10'hd5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_213; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2355 = 10'hd6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_214; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2356 = 10'hd7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_215; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2357 = 10'hd8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_216; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2358 = 10'hd9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_217; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2359 = 10'hda == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_218; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2360 = 10'hdb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_219; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2361 = 10'hdc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_220; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2362 = 10'hdd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_221; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2363 = 10'hde == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_222; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2364 = 10'hdf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_223; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2365 = 10'he0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_224; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2366 = 10'he1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_225; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2367 = 10'he2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_226; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2368 = 10'he3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_227; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2369 = 10'he4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_228; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2370 = 10'he5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_229; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2371 = 10'he6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_230; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2372 = 10'he7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_231; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2373 = 10'he8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_232; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2374 = 10'he9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_233; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2375 = 10'hea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_234; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2376 = 10'heb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_235; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2377 = 10'hec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_236; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2378 = 10'hed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_237; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2379 = 10'hee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_238; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2380 = 10'hef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_239; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2381 = 10'hf0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_240; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2382 = 10'hf1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_241; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2383 = 10'hf2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_242; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2384 = 10'hf3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_243; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2385 = 10'hf4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_244; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2386 = 10'hf5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_245; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2387 = 10'hf6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_246; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2388 = 10'hf7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_247; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2389 = 10'hf8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_248; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2390 = 10'hf9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_249; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2391 = 10'hfa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_250; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2392 = 10'hfb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_251; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2393 = 10'hfc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_252; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2394 = 10'hfd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_253; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2395 = 10'hfe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_254; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2396 = 10'hff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_255; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2397 = 10'h100 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_256; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2398 = 10'h101 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_257; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2399 = 10'h102 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_258; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2400 = 10'h103 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_259; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2401 = 10'h104 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_260; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2402 = 10'h105 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_261; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2403 = 10'h106 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_262; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2404 = 10'h107 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_263; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2405 = 10'h108 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_264; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2406 = 10'h109 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_265; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2407 = 10'h10a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_266; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2408 = 10'h10b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_267; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2409 = 10'h10c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_268; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2410 = 10'h10d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_269; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2411 = 10'h10e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_270; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2412 = 10'h10f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_271; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2413 = 10'h110 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_272; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2414 = 10'h111 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_273; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2415 = 10'h112 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_274; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2416 = 10'h113 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_275; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2417 = 10'h114 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_276; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2418 = 10'h115 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_277; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2419 = 10'h116 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_278; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2420 = 10'h117 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_279; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2421 = 10'h118 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_280; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2422 = 10'h119 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_281; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2423 = 10'h11a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_282; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2424 = 10'h11b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_283; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2425 = 10'h11c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_284; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2426 = 10'h11d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_285; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2427 = 10'h11e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_286; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2428 = 10'h11f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_287; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2429 = 10'h120 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_288; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2430 = 10'h121 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_289; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2431 = 10'h122 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_290; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2432 = 10'h123 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_291; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2433 = 10'h124 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_292; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2434 = 10'h125 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_293; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2435 = 10'h126 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_294; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2436 = 10'h127 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_295; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2437 = 10'h128 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_296; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2438 = 10'h129 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_297; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2439 = 10'h12a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_298; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2440 = 10'h12b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_299; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2441 = 10'h12c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_300; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2442 = 10'h12d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_301; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2443 = 10'h12e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_302; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2444 = 10'h12f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_303; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2445 = 10'h130 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_304; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2446 = 10'h131 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_305; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2447 = 10'h132 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_306; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2448 = 10'h133 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_307; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2449 = 10'h134 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_308; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2450 = 10'h135 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_309; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2451 = 10'h136 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_310; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2452 = 10'h137 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_311; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2453 = 10'h138 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_312; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2454 = 10'h139 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_313; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2455 = 10'h13a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_314; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2456 = 10'h13b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_315; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2457 = 10'h13c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_316; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2458 = 10'h13d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_317; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2459 = 10'h13e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_318; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2460 = 10'h13f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_319; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2461 = 10'h140 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_320; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2462 = 10'h141 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_321; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2463 = 10'h142 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_322; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2464 = 10'h143 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_323; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2465 = 10'h144 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_324; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2466 = 10'h145 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_325; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2467 = 10'h146 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_326; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2468 = 10'h147 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_327; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2469 = 10'h148 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_328; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2470 = 10'h149 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_329; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2471 = 10'h14a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_330; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2472 = 10'h14b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_331; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2473 = 10'h14c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_332; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2474 = 10'h14d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_333; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2475 = 10'h14e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_334; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2476 = 10'h14f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_335; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2477 = 10'h150 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_336; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2478 = 10'h151 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_337; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2479 = 10'h152 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_338; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2480 = 10'h153 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_339; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2481 = 10'h154 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_340; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2482 = 10'h155 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_341; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2483 = 10'h156 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_342; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2484 = 10'h157 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_343; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2485 = 10'h158 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_344; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2486 = 10'h159 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_345; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2487 = 10'h15a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_346; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2488 = 10'h15b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_347; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2489 = 10'h15c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_348; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2490 = 10'h15d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_349; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2491 = 10'h15e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_350; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2492 = 10'h15f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_351; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2493 = 10'h160 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_352; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2494 = 10'h161 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_353; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2495 = 10'h162 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_354; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2496 = 10'h163 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_355; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2497 = 10'h164 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_356; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2498 = 10'h165 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_357; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2499 = 10'h166 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_358; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2500 = 10'h167 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_359; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2501 = 10'h168 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_360; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2502 = 10'h169 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_361; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2503 = 10'h16a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_362; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2504 = 10'h16b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_363; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2505 = 10'h16c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_364; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2506 = 10'h16d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_365; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2507 = 10'h16e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_366; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2508 = 10'h16f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_367; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2509 = 10'h170 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_368; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2510 = 10'h171 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_369; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2511 = 10'h172 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_370; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2512 = 10'h173 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_371; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2513 = 10'h174 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_372; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2514 = 10'h175 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_373; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2515 = 10'h176 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_374; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2516 = 10'h177 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_375; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2517 = 10'h178 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_376; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2518 = 10'h179 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_377; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2519 = 10'h17a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_378; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2520 = 10'h17b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_379; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2521 = 10'h17c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_380; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2522 = 10'h17d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_381; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2523 = 10'h17e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_382; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2524 = 10'h17f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_383; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2525 = 10'h180 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_384; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2526 = 10'h181 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_385; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2527 = 10'h182 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_386; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2528 = 10'h183 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_387; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2529 = 10'h184 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_388; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2530 = 10'h185 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_389; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2531 = 10'h186 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_390; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2532 = 10'h187 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_391; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2533 = 10'h188 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_392; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2534 = 10'h189 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_393; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2535 = 10'h18a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_394; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2536 = 10'h18b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_395; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2537 = 10'h18c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_396; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2538 = 10'h18d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_397; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2539 = 10'h18e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_398; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2540 = 10'h18f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_399; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2541 = 10'h190 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_400; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2542 = 10'h191 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_401; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2543 = 10'h192 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_402; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2544 = 10'h193 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_403; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2545 = 10'h194 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_404; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2546 = 10'h195 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_405; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2547 = 10'h196 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_406; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2548 = 10'h197 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_407; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2549 = 10'h198 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_408; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2550 = 10'h199 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_409; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2551 = 10'h19a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_410; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2552 = 10'h19b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_411; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2553 = 10'h19c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_412; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2554 = 10'h19d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_413; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2555 = 10'h19e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_414; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2556 = 10'h19f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_415; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2557 = 10'h1a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_416; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2558 = 10'h1a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_417; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2559 = 10'h1a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_418; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2560 = 10'h1a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_419; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2561 = 10'h1a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_420; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2562 = 10'h1a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_421; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2563 = 10'h1a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_422; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2564 = 10'h1a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_423; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2565 = 10'h1a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_424; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2566 = 10'h1a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_425; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2567 = 10'h1aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_426; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2568 = 10'h1ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_427; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2569 = 10'h1ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_428; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2570 = 10'h1ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_429; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2571 = 10'h1ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_430; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2572 = 10'h1af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_431; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2573 = 10'h1b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_432; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2574 = 10'h1b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_433; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2575 = 10'h1b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_434; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2576 = 10'h1b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_435; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2577 = 10'h1b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_436; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2578 = 10'h1b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_437; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2579 = 10'h1b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_438; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2580 = 10'h1b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_439; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2581 = 10'h1b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_440; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2582 = 10'h1b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_441; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2583 = 10'h1ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_442; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2584 = 10'h1bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_443; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2585 = 10'h1bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_444; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2586 = 10'h1bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_445; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2587 = 10'h1be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_446; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2588 = 10'h1bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_447; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2589 = 10'h1c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_448; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2590 = 10'h1c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_449; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2591 = 10'h1c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_450; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2592 = 10'h1c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_451; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2593 = 10'h1c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_452; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2594 = 10'h1c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_453; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2595 = 10'h1c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_454; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2596 = 10'h1c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_455; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2597 = 10'h1c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_456; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2598 = 10'h1c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_457; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2599 = 10'h1ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_458; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2600 = 10'h1cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_459; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2601 = 10'h1cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_460; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2602 = 10'h1cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_461; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2603 = 10'h1ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_462; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2604 = 10'h1cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_463; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2605 = 10'h1d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_464; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2606 = 10'h1d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_465; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2607 = 10'h1d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_466; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2608 = 10'h1d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_467; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2609 = 10'h1d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_468; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2610 = 10'h1d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_469; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2611 = 10'h1d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_470; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2612 = 10'h1d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_471; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2613 = 10'h1d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_472; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2614 = 10'h1d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_473; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2615 = 10'h1da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_474; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2616 = 10'h1db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_475; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2617 = 10'h1dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_476; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2618 = 10'h1dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_477; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2619 = 10'h1de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_478; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2620 = 10'h1df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_479; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2621 = 10'h1e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_480; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2622 = 10'h1e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_481; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2623 = 10'h1e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_482; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2624 = 10'h1e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_483; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2625 = 10'h1e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_484; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2626 = 10'h1e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_485; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2627 = 10'h1e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_486; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2628 = 10'h1e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_487; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2629 = 10'h1e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_488; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2630 = 10'h1e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_489; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2631 = 10'h1ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_490; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2632 = 10'h1eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_491; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2633 = 10'h1ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_492; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2634 = 10'h1ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_493; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2635 = 10'h1ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_494; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2636 = 10'h1ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_495; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2637 = 10'h1f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_496; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2638 = 10'h1f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_497; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2639 = 10'h1f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_498; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2640 = 10'h1f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_499; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2641 = 10'h1f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_500; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2642 = 10'h1f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_501; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2643 = 10'h1f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_502; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2644 = 10'h1f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_503; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2645 = 10'h1f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_504; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2646 = 10'h1f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_505; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2647 = 10'h1fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_506; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2648 = 10'h1fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_507; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2649 = 10'h1fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_508; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2650 = 10'h1fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_509; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2651 = 10'h1fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_510; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2652 = 10'h1ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_511; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2653 = 10'h200 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_512; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2654 = 10'h201 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_513; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2655 = 10'h202 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_514; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2656 = 10'h203 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_515; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2657 = 10'h204 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_516; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2658 = 10'h205 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_517; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2659 = 10'h206 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_518; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2660 = 10'h207 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_519; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2661 = 10'h208 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_520; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2662 = 10'h209 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_521; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2663 = 10'h20a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_522; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2664 = 10'h20b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_523; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2665 = 10'h20c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_524; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2666 = 10'h20d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_525; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2667 = 10'h20e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_526; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2668 = 10'h20f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_527; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2669 = 10'h210 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_528; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2670 = 10'h211 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_529; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2671 = 10'h212 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_530; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2672 = 10'h213 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_531; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2673 = 10'h214 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_532; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2674 = 10'h215 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_533; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2675 = 10'h216 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_534; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2676 = 10'h217 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_535; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2677 = 10'h218 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_536; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2678 = 10'h219 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_537; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2679 = 10'h21a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_538; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2680 = 10'h21b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_539; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2681 = 10'h21c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_540; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2682 = 10'h21d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_541; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2683 = 10'h21e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_542; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2684 = 10'h21f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_543; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2685 = 10'h220 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_544; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2686 = 10'h221 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_545; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2687 = 10'h222 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_546; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2688 = 10'h223 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_547; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2689 = 10'h224 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_548; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2690 = 10'h225 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_549; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2691 = 10'h226 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_550; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2692 = 10'h227 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_551; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2693 = 10'h228 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_552; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2694 = 10'h229 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_553; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2695 = 10'h22a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_554; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2696 = 10'h22b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_555; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2697 = 10'h22c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_556; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2698 = 10'h22d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_557; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2699 = 10'h22e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_558; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2700 = 10'h22f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_559; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2701 = 10'h230 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_560; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2702 = 10'h231 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_561; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2703 = 10'h232 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_562; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2704 = 10'h233 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_563; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2705 = 10'h234 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_564; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2706 = 10'h235 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_565; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2707 = 10'h236 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_566; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2708 = 10'h237 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_567; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2709 = 10'h238 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_568; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2710 = 10'h239 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_569; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2711 = 10'h23a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_570; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2712 = 10'h23b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_571; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2713 = 10'h23c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_572; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2714 = 10'h23d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_573; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2715 = 10'h23e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_574; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2716 = 10'h23f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_575; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2717 = 10'h240 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_576; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2718 = 10'h241 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_577; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2719 = 10'h242 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_578; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2720 = 10'h243 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_579; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2721 = 10'h244 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_580; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2722 = 10'h245 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_581; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2723 = 10'h246 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_582; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2724 = 10'h247 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_583; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2725 = 10'h248 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_584; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2726 = 10'h249 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_585; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2727 = 10'h24a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_586; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2728 = 10'h24b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_587; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2729 = 10'h24c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_588; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2730 = 10'h24d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_589; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2731 = 10'h24e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_590; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2732 = 10'h24f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_591; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2733 = 10'h250 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_592; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2734 = 10'h251 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_593; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2735 = 10'h252 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_594; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2736 = 10'h253 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_595; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2737 = 10'h254 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_596; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2738 = 10'h255 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_597; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2739 = 10'h256 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_598; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2740 = 10'h257 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_599; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2741 = 10'h258 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_600; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2742 = 10'h259 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_601; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2743 = 10'h25a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_602; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2744 = 10'h25b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_603; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2745 = 10'h25c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_604; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2746 = 10'h25d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_605; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2747 = 10'h25e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_606; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2748 = 10'h25f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_607; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2749 = 10'h260 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_608; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2750 = 10'h261 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_609; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2751 = 10'h262 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_610; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2752 = 10'h263 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_611; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2753 = 10'h264 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_612; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2754 = 10'h265 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_613; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2755 = 10'h266 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_614; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2756 = 10'h267 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_615; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2757 = 10'h268 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_616; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2758 = 10'h269 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_617; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2759 = 10'h26a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_618; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2760 = 10'h26b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_619; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2761 = 10'h26c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_620; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2762 = 10'h26d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_621; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2763 = 10'h26e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_622; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2764 = 10'h26f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_623; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2765 = 10'h270 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_624; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2766 = 10'h271 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_625; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2767 = 10'h272 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_626; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2768 = 10'h273 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_627; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2769 = 10'h274 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_628; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2770 = 10'h275 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_629; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2771 = 10'h276 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_630; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2772 = 10'h277 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_631; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2773 = 10'h278 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_632; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2774 = 10'h279 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_633; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2775 = 10'h27a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_634; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2776 = 10'h27b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_635; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2777 = 10'h27c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_636; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2778 = 10'h27d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_637; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2779 = 10'h27e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_638; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2780 = 10'h27f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_639; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2781 = 10'h280 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_640; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2782 = 10'h281 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_641; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2783 = 10'h282 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_642; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2784 = 10'h283 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_643; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2785 = 10'h284 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_644; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2786 = 10'h285 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_645; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2787 = 10'h286 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_646; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2788 = 10'h287 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_647; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2789 = 10'h288 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_648; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2790 = 10'h289 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_649; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2791 = 10'h28a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_650; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2792 = 10'h28b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_651; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2793 = 10'h28c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_652; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2794 = 10'h28d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_653; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2795 = 10'h28e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_654; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2796 = 10'h28f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_655; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2797 = 10'h290 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_656; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2798 = 10'h291 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_657; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2799 = 10'h292 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_658; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2800 = 10'h293 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_659; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2801 = 10'h294 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_660; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2802 = 10'h295 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_661; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2803 = 10'h296 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_662; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2804 = 10'h297 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_663; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2805 = 10'h298 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_664; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2806 = 10'h299 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_665; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2807 = 10'h29a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_666; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2808 = 10'h29b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_667; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2809 = 10'h29c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_668; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2810 = 10'h29d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_669; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2811 = 10'h29e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_670; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2812 = 10'h29f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_671; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2813 = 10'h2a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_672; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2814 = 10'h2a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_673; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2815 = 10'h2a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_674; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2816 = 10'h2a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_675; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2817 = 10'h2a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_676; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2818 = 10'h2a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_677; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2819 = 10'h2a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_678; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2820 = 10'h2a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_679; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2821 = 10'h2a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_680; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2822 = 10'h2a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_681; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2823 = 10'h2aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_682; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2824 = 10'h2ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_683; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2825 = 10'h2ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_684; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2826 = 10'h2ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_685; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2827 = 10'h2ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_686; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2828 = 10'h2af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_687; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2829 = 10'h2b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_688; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2830 = 10'h2b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_689; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2831 = 10'h2b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_690; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2832 = 10'h2b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_691; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2833 = 10'h2b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_692; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2834 = 10'h2b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_693; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2835 = 10'h2b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_694; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2836 = 10'h2b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_695; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2837 = 10'h2b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_696; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2838 = 10'h2b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_697; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2839 = 10'h2ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_698; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2840 = 10'h2bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_699; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2841 = 10'h2bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_700; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2842 = 10'h2bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_701; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2843 = 10'h2be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_702; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2844 = 10'h2bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_703; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2845 = 10'h2c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_704; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2846 = 10'h2c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_705; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2847 = 10'h2c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_706; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2848 = 10'h2c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_707; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2849 = 10'h2c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_708; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2850 = 10'h2c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_709; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2851 = 10'h2c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_710; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2852 = 10'h2c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_711; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2853 = 10'h2c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_712; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2854 = 10'h2c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_713; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2855 = 10'h2ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_714; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2856 = 10'h2cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_715; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2857 = 10'h2cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_716; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2858 = 10'h2cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_717; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2859 = 10'h2ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_718; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2860 = 10'h2cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_719; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2861 = 10'h2d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_720; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2862 = 10'h2d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_721; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2863 = 10'h2d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_722; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2864 = 10'h2d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_723; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2865 = 10'h2d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_724; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2866 = 10'h2d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_725; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2867 = 10'h2d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_726; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2868 = 10'h2d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_727; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2869 = 10'h2d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_728; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2870 = 10'h2d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_729; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2871 = 10'h2da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_730; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2872 = 10'h2db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_731; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2873 = 10'h2dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_732; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2874 = 10'h2dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_733; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2875 = 10'h2de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_734; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2876 = 10'h2df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_735; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2877 = 10'h2e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_736; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2878 = 10'h2e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_737; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2879 = 10'h2e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_738; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2880 = 10'h2e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_739; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2881 = 10'h2e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_740; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2882 = 10'h2e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_741; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2883 = 10'h2e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_742; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2884 = 10'h2e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_743; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2885 = 10'h2e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_744; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2886 = 10'h2e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_745; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2887 = 10'h2ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_746; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2888 = 10'h2eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_747; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2889 = 10'h2ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_748; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2890 = 10'h2ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_749; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2891 = 10'h2ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_750; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2892 = 10'h2ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_751; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2893 = 10'h2f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_752; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2894 = 10'h2f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_753; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2895 = 10'h2f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_754; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2896 = 10'h2f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_755; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2897 = 10'h2f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_756; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2898 = 10'h2f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_757; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2899 = 10'h2f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_758; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2900 = 10'h2f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_759; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2901 = 10'h2f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_760; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2902 = 10'h2f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_761; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2903 = 10'h2fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_762; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2904 = 10'h2fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_763; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2905 = 10'h2fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_764; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2906 = 10'h2fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_765; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2907 = 10'h2fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_766; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2908 = 10'h2ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_767; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2909 = 10'h300 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_768; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2910 = 10'h301 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_769; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2911 = 10'h302 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_770; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2912 = 10'h303 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_771; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2913 = 10'h304 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_772; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2914 = 10'h305 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_773; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2915 = 10'h306 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_774; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2916 = 10'h307 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_775; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2917 = 10'h308 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_776; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2918 = 10'h309 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_777; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2919 = 10'h30a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_778; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2920 = 10'h30b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_779; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2921 = 10'h30c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_780; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2922 = 10'h30d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_781; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2923 = 10'h30e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_782; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2924 = 10'h30f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_783; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2925 = 10'h310 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_784; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2926 = 10'h311 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_785; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2927 = 10'h312 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_786; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2928 = 10'h313 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_787; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2929 = 10'h314 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_788; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2930 = 10'h315 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_789; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2931 = 10'h316 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_790; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2932 = 10'h317 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_791; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2933 = 10'h318 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_792; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2934 = 10'h319 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_793; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2935 = 10'h31a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_794; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2936 = 10'h31b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_795; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2937 = 10'h31c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_796; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2938 = 10'h31d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_797; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2939 = 10'h31e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_798; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2940 = 10'h31f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_799; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2941 = 10'h320 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_800; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2942 = 10'h321 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_801; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2943 = 10'h322 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_802; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2944 = 10'h323 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_803; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2945 = 10'h324 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_804; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2946 = 10'h325 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_805; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2947 = 10'h326 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_806; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2948 = 10'h327 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_807; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2949 = 10'h328 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_808; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2950 = 10'h329 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_809; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2951 = 10'h32a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_810; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2952 = 10'h32b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_811; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2953 = 10'h32c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_812; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2954 = 10'h32d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_813; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2955 = 10'h32e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_814; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2956 = 10'h32f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_815; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2957 = 10'h330 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_816; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2958 = 10'h331 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_817; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2959 = 10'h332 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_818; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2960 = 10'h333 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_819; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2961 = 10'h334 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_820; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2962 = 10'h335 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_821; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2963 = 10'h336 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_822; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2964 = 10'h337 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_823; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2965 = 10'h338 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_824; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2966 = 10'h339 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_825; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2967 = 10'h33a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_826; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2968 = 10'h33b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_827; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2969 = 10'h33c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_828; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2970 = 10'h33d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_829; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2971 = 10'h33e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_830; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2972 = 10'h33f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_831; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2973 = 10'h340 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_832; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2974 = 10'h341 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_833; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2975 = 10'h342 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_834; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2976 = 10'h343 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_835; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2977 = 10'h344 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_836; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2978 = 10'h345 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_837; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2979 = 10'h346 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_838; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2980 = 10'h347 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_839; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2981 = 10'h348 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_840; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2982 = 10'h349 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_841; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2983 = 10'h34a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_842; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2984 = 10'h34b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_843; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2985 = 10'h34c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_844; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2986 = 10'h34d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_845; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2987 = 10'h34e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_846; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2988 = 10'h34f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_847; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2989 = 10'h350 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_848; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2990 = 10'h351 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_849; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2991 = 10'h352 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_850; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2992 = 10'h353 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_851; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2993 = 10'h354 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_852; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2994 = 10'h355 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_853; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2995 = 10'h356 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_854; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2996 = 10'h357 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_855; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2997 = 10'h358 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_856; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2998 = 10'h359 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_857; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_2999 = 10'h35a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_858; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3000 = 10'h35b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_859; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3001 = 10'h35c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_860; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3002 = 10'h35d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_861; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3003 = 10'h35e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_862; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3004 = 10'h35f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_863; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3005 = 10'h360 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_864; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3006 = 10'h361 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_865; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3007 = 10'h362 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_866; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3008 = 10'h363 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_867; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3009 = 10'h364 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_868; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3010 = 10'h365 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_869; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3011 = 10'h366 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_870; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3012 = 10'h367 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_871; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3013 = 10'h368 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_872; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3014 = 10'h369 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_873; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3015 = 10'h36a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_874; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3016 = 10'h36b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_875; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3017 = 10'h36c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_876; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3018 = 10'h36d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_877; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3019 = 10'h36e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_878; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3020 = 10'h36f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_879; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3021 = 10'h370 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_880; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3022 = 10'h371 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_881; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3023 = 10'h372 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_882; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3024 = 10'h373 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_883; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3025 = 10'h374 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_884; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3026 = 10'h375 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_885; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3027 = 10'h376 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_886; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3028 = 10'h377 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_887; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3029 = 10'h378 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_888; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3030 = 10'h379 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_889; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3031 = 10'h37a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_890; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3032 = 10'h37b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_891; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3033 = 10'h37c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_892; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3034 = 10'h37d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_893; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3035 = 10'h37e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_894; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3036 = 10'h37f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_895; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3037 = 10'h380 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_896; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3038 = 10'h381 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_897; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3039 = 10'h382 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_898; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3040 = 10'h383 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_899; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3041 = 10'h384 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_900; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3042 = 10'h385 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_901; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3043 = 10'h386 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_902; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3044 = 10'h387 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_903; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3045 = 10'h388 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_904; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3046 = 10'h389 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_905; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3047 = 10'h38a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_906; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3048 = 10'h38b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_907; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3049 = 10'h38c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_908; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3050 = 10'h38d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_909; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3051 = 10'h38e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_910; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3052 = 10'h38f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_911; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3053 = 10'h390 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_912; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3054 = 10'h391 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_913; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3055 = 10'h392 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_914; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3056 = 10'h393 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_915; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3057 = 10'h394 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_916; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3058 = 10'h395 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_917; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3059 = 10'h396 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_918; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3060 = 10'h397 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_919; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3061 = 10'h398 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_920; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3062 = 10'h399 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_921; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3063 = 10'h39a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_922; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3064 = 10'h39b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_923; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3065 = 10'h39c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_924; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3066 = 10'h39d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_925; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3067 = 10'h39e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_926; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3068 = 10'h39f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_927; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3069 = 10'h3a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_928; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3070 = 10'h3a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_929; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3071 = 10'h3a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_930; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3072 = 10'h3a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_931; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3073 = 10'h3a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_932; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3074 = 10'h3a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_933; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3075 = 10'h3a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_934; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3076 = 10'h3a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_935; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3077 = 10'h3a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_936; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3078 = 10'h3a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_937; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3079 = 10'h3aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_938; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3080 = 10'h3ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_939; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3081 = 10'h3ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_940; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3082 = 10'h3ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_941; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3083 = 10'h3ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_942; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3084 = 10'h3af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_943; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3085 = 10'h3b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_944; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3086 = 10'h3b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_945; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3087 = 10'h3b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_946; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3088 = 10'h3b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_947; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3089 = 10'h3b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_948; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3090 = 10'h3b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_949; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3091 = 10'h3b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_950; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3092 = 10'h3b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_951; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3093 = 10'h3b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_952; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3094 = 10'h3b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_953; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3095 = 10'h3ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_954; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3096 = 10'h3bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_955; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3097 = 10'h3bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_956; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3098 = 10'h3bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_957; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3099 = 10'h3be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_958; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3100 = 10'h3bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_959; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3101 = 10'h3c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_960; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3102 = 10'h3c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_961; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3103 = 10'h3c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_962; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3104 = 10'h3c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_963; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3105 = 10'h3c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_964; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3106 = 10'h3c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_965; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3107 = 10'h3c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_966; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3108 = 10'h3c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_967; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3109 = 10'h3c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_968; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3110 = 10'h3c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_969; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3111 = 10'h3ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_970; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3112 = 10'h3cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_971; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3113 = 10'h3cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_972; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3114 = 10'h3cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_973; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3115 = 10'h3ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_974; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3116 = 10'h3cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_975; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3117 = 10'h3d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_976; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3118 = 10'h3d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_977; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3119 = 10'h3d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_978; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3120 = 10'h3d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_979; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3121 = 10'h3d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_980; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3122 = 10'h3d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_981; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3123 = 10'h3d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_982; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3124 = 10'h3d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_983; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3125 = 10'h3d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_984; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3126 = 10'h3d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_985; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3127 = 10'h3da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_986; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3128 = 10'h3db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_987; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3129 = 10'h3dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_988; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3130 = 10'h3dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_989; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3131 = 10'h3de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_990; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3132 = 10'h3df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_991; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3133 = 10'h3e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_992; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3134 = 10'h3e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_993; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3135 = 10'h3e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_994; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3136 = 10'h3e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_995; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3137 = 10'h3e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_996; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3138 = 10'h3e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_997; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3139 = 10'h3e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_998; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3140 = 10'h3e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_999; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3141 = 10'h3e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1000; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3142 = 10'h3e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1001; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3143 = 10'h3ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1002; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3144 = 10'h3eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1003; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3145 = 10'h3ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1004; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3146 = 10'h3ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1005; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3147 = 10'h3ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1006; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3148 = 10'h3ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1007; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3149 = 10'h3f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1008; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3150 = 10'h3f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1009; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3151 = 10'h3f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1010; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3152 = 10'h3f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1011; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3153 = 10'h3f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1012; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3154 = 10'h3f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1013; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3155 = 10'h3f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1014; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3156 = 10'h3f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1015; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3157 = 10'h3f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1016; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3158 = 10'h3f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1017; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3159 = 10'h3fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1018; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3160 = 10'h3fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1019; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3161 = 10'h3fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1020; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3162 = 10'h3fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1021; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3163 = 10'h3fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1022; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3164 = 10'h3ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1023; // @[cpu.scala 221:{37,37} 69:24]
  wire [31:0] _GEN_3165 = EXMEMop == 7'h23 ? _GEN_2141 : DMemory_0; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3166 = EXMEMop == 7'h23 ? _GEN_2142 : DMemory_1; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3167 = EXMEMop == 7'h23 ? _GEN_2143 : DMemory_2; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3168 = EXMEMop == 7'h23 ? _GEN_2144 : DMemory_3; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3169 = EXMEMop == 7'h23 ? _GEN_2145 : DMemory_4; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3170 = EXMEMop == 7'h23 ? _GEN_2146 : DMemory_5; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3171 = EXMEMop == 7'h23 ? _GEN_2147 : DMemory_6; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3172 = EXMEMop == 7'h23 ? _GEN_2148 : DMemory_7; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3173 = EXMEMop == 7'h23 ? _GEN_2149 : DMemory_8; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3174 = EXMEMop == 7'h23 ? _GEN_2150 : DMemory_9; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3175 = EXMEMop == 7'h23 ? _GEN_2151 : DMemory_10; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3176 = EXMEMop == 7'h23 ? _GEN_2152 : DMemory_11; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3177 = EXMEMop == 7'h23 ? _GEN_2153 : DMemory_12; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3178 = EXMEMop == 7'h23 ? _GEN_2154 : DMemory_13; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3179 = EXMEMop == 7'h23 ? _GEN_2155 : DMemory_14; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3180 = EXMEMop == 7'h23 ? _GEN_2156 : DMemory_15; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3181 = EXMEMop == 7'h23 ? _GEN_2157 : DMemory_16; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3182 = EXMEMop == 7'h23 ? _GEN_2158 : DMemory_17; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3183 = EXMEMop == 7'h23 ? _GEN_2159 : DMemory_18; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3184 = EXMEMop == 7'h23 ? _GEN_2160 : DMemory_19; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3185 = EXMEMop == 7'h23 ? _GEN_2161 : DMemory_20; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3186 = EXMEMop == 7'h23 ? _GEN_2162 : DMemory_21; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3187 = EXMEMop == 7'h23 ? _GEN_2163 : DMemory_22; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3188 = EXMEMop == 7'h23 ? _GEN_2164 : DMemory_23; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3189 = EXMEMop == 7'h23 ? _GEN_2165 : DMemory_24; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3190 = EXMEMop == 7'h23 ? _GEN_2166 : DMemory_25; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3191 = EXMEMop == 7'h23 ? _GEN_2167 : DMemory_26; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3192 = EXMEMop == 7'h23 ? _GEN_2168 : DMemory_27; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3193 = EXMEMop == 7'h23 ? _GEN_2169 : DMemory_28; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3194 = EXMEMop == 7'h23 ? _GEN_2170 : DMemory_29; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3195 = EXMEMop == 7'h23 ? _GEN_2171 : DMemory_30; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3196 = EXMEMop == 7'h23 ? _GEN_2172 : DMemory_31; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3197 = EXMEMop == 7'h23 ? _GEN_2173 : DMemory_32; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3198 = EXMEMop == 7'h23 ? _GEN_2174 : DMemory_33; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3199 = EXMEMop == 7'h23 ? _GEN_2175 : DMemory_34; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3200 = EXMEMop == 7'h23 ? _GEN_2176 : DMemory_35; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3201 = EXMEMop == 7'h23 ? _GEN_2177 : DMemory_36; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3202 = EXMEMop == 7'h23 ? _GEN_2178 : DMemory_37; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3203 = EXMEMop == 7'h23 ? _GEN_2179 : DMemory_38; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3204 = EXMEMop == 7'h23 ? _GEN_2180 : DMemory_39; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3205 = EXMEMop == 7'h23 ? _GEN_2181 : DMemory_40; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3206 = EXMEMop == 7'h23 ? _GEN_2182 : DMemory_41; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3207 = EXMEMop == 7'h23 ? _GEN_2183 : DMemory_42; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3208 = EXMEMop == 7'h23 ? _GEN_2184 : DMemory_43; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3209 = EXMEMop == 7'h23 ? _GEN_2185 : DMemory_44; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3210 = EXMEMop == 7'h23 ? _GEN_2186 : DMemory_45; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3211 = EXMEMop == 7'h23 ? _GEN_2187 : DMemory_46; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3212 = EXMEMop == 7'h23 ? _GEN_2188 : DMemory_47; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3213 = EXMEMop == 7'h23 ? _GEN_2189 : DMemory_48; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3214 = EXMEMop == 7'h23 ? _GEN_2190 : DMemory_49; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3215 = EXMEMop == 7'h23 ? _GEN_2191 : DMemory_50; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3216 = EXMEMop == 7'h23 ? _GEN_2192 : DMemory_51; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3217 = EXMEMop == 7'h23 ? _GEN_2193 : DMemory_52; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3218 = EXMEMop == 7'h23 ? _GEN_2194 : DMemory_53; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3219 = EXMEMop == 7'h23 ? _GEN_2195 : DMemory_54; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3220 = EXMEMop == 7'h23 ? _GEN_2196 : DMemory_55; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3221 = EXMEMop == 7'h23 ? _GEN_2197 : DMemory_56; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3222 = EXMEMop == 7'h23 ? _GEN_2198 : DMemory_57; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3223 = EXMEMop == 7'h23 ? _GEN_2199 : DMemory_58; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3224 = EXMEMop == 7'h23 ? _GEN_2200 : DMemory_59; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3225 = EXMEMop == 7'h23 ? _GEN_2201 : DMemory_60; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3226 = EXMEMop == 7'h23 ? _GEN_2202 : DMemory_61; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3227 = EXMEMop == 7'h23 ? _GEN_2203 : DMemory_62; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3228 = EXMEMop == 7'h23 ? _GEN_2204 : DMemory_63; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3229 = EXMEMop == 7'h23 ? _GEN_2205 : DMemory_64; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3230 = EXMEMop == 7'h23 ? _GEN_2206 : DMemory_65; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3231 = EXMEMop == 7'h23 ? _GEN_2207 : DMemory_66; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3232 = EXMEMop == 7'h23 ? _GEN_2208 : DMemory_67; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3233 = EXMEMop == 7'h23 ? _GEN_2209 : DMemory_68; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3234 = EXMEMop == 7'h23 ? _GEN_2210 : DMemory_69; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3235 = EXMEMop == 7'h23 ? _GEN_2211 : DMemory_70; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3236 = EXMEMop == 7'h23 ? _GEN_2212 : DMemory_71; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3237 = EXMEMop == 7'h23 ? _GEN_2213 : DMemory_72; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3238 = EXMEMop == 7'h23 ? _GEN_2214 : DMemory_73; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3239 = EXMEMop == 7'h23 ? _GEN_2215 : DMemory_74; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3240 = EXMEMop == 7'h23 ? _GEN_2216 : DMemory_75; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3241 = EXMEMop == 7'h23 ? _GEN_2217 : DMemory_76; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3242 = EXMEMop == 7'h23 ? _GEN_2218 : DMemory_77; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3243 = EXMEMop == 7'h23 ? _GEN_2219 : DMemory_78; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3244 = EXMEMop == 7'h23 ? _GEN_2220 : DMemory_79; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3245 = EXMEMop == 7'h23 ? _GEN_2221 : DMemory_80; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3246 = EXMEMop == 7'h23 ? _GEN_2222 : DMemory_81; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3247 = EXMEMop == 7'h23 ? _GEN_2223 : DMemory_82; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3248 = EXMEMop == 7'h23 ? _GEN_2224 : DMemory_83; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3249 = EXMEMop == 7'h23 ? _GEN_2225 : DMemory_84; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3250 = EXMEMop == 7'h23 ? _GEN_2226 : DMemory_85; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3251 = EXMEMop == 7'h23 ? _GEN_2227 : DMemory_86; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3252 = EXMEMop == 7'h23 ? _GEN_2228 : DMemory_87; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3253 = EXMEMop == 7'h23 ? _GEN_2229 : DMemory_88; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3254 = EXMEMop == 7'h23 ? _GEN_2230 : DMemory_89; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3255 = EXMEMop == 7'h23 ? _GEN_2231 : DMemory_90; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3256 = EXMEMop == 7'h23 ? _GEN_2232 : DMemory_91; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3257 = EXMEMop == 7'h23 ? _GEN_2233 : DMemory_92; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3258 = EXMEMop == 7'h23 ? _GEN_2234 : DMemory_93; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3259 = EXMEMop == 7'h23 ? _GEN_2235 : DMemory_94; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3260 = EXMEMop == 7'h23 ? _GEN_2236 : DMemory_95; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3261 = EXMEMop == 7'h23 ? _GEN_2237 : DMemory_96; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3262 = EXMEMop == 7'h23 ? _GEN_2238 : DMemory_97; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3263 = EXMEMop == 7'h23 ? _GEN_2239 : DMemory_98; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3264 = EXMEMop == 7'h23 ? _GEN_2240 : DMemory_99; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3265 = EXMEMop == 7'h23 ? _GEN_2241 : DMemory_100; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3266 = EXMEMop == 7'h23 ? _GEN_2242 : DMemory_101; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3267 = EXMEMop == 7'h23 ? _GEN_2243 : DMemory_102; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3268 = EXMEMop == 7'h23 ? _GEN_2244 : DMemory_103; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3269 = EXMEMop == 7'h23 ? _GEN_2245 : DMemory_104; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3270 = EXMEMop == 7'h23 ? _GEN_2246 : DMemory_105; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3271 = EXMEMop == 7'h23 ? _GEN_2247 : DMemory_106; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3272 = EXMEMop == 7'h23 ? _GEN_2248 : DMemory_107; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3273 = EXMEMop == 7'h23 ? _GEN_2249 : DMemory_108; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3274 = EXMEMop == 7'h23 ? _GEN_2250 : DMemory_109; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3275 = EXMEMop == 7'h23 ? _GEN_2251 : DMemory_110; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3276 = EXMEMop == 7'h23 ? _GEN_2252 : DMemory_111; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3277 = EXMEMop == 7'h23 ? _GEN_2253 : DMemory_112; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3278 = EXMEMop == 7'h23 ? _GEN_2254 : DMemory_113; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3279 = EXMEMop == 7'h23 ? _GEN_2255 : DMemory_114; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3280 = EXMEMop == 7'h23 ? _GEN_2256 : DMemory_115; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3281 = EXMEMop == 7'h23 ? _GEN_2257 : DMemory_116; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3282 = EXMEMop == 7'h23 ? _GEN_2258 : DMemory_117; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3283 = EXMEMop == 7'h23 ? _GEN_2259 : DMemory_118; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3284 = EXMEMop == 7'h23 ? _GEN_2260 : DMemory_119; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3285 = EXMEMop == 7'h23 ? _GEN_2261 : DMemory_120; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3286 = EXMEMop == 7'h23 ? _GEN_2262 : DMemory_121; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3287 = EXMEMop == 7'h23 ? _GEN_2263 : DMemory_122; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3288 = EXMEMop == 7'h23 ? _GEN_2264 : DMemory_123; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3289 = EXMEMop == 7'h23 ? _GEN_2265 : DMemory_124; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3290 = EXMEMop == 7'h23 ? _GEN_2266 : DMemory_125; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3291 = EXMEMop == 7'h23 ? _GEN_2267 : DMemory_126; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3292 = EXMEMop == 7'h23 ? _GEN_2268 : DMemory_127; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3293 = EXMEMop == 7'h23 ? _GEN_2269 : DMemory_128; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3294 = EXMEMop == 7'h23 ? _GEN_2270 : DMemory_129; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3295 = EXMEMop == 7'h23 ? _GEN_2271 : DMemory_130; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3296 = EXMEMop == 7'h23 ? _GEN_2272 : DMemory_131; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3297 = EXMEMop == 7'h23 ? _GEN_2273 : DMemory_132; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3298 = EXMEMop == 7'h23 ? _GEN_2274 : DMemory_133; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3299 = EXMEMop == 7'h23 ? _GEN_2275 : DMemory_134; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3300 = EXMEMop == 7'h23 ? _GEN_2276 : DMemory_135; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3301 = EXMEMop == 7'h23 ? _GEN_2277 : DMemory_136; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3302 = EXMEMop == 7'h23 ? _GEN_2278 : DMemory_137; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3303 = EXMEMop == 7'h23 ? _GEN_2279 : DMemory_138; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3304 = EXMEMop == 7'h23 ? _GEN_2280 : DMemory_139; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3305 = EXMEMop == 7'h23 ? _GEN_2281 : DMemory_140; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3306 = EXMEMop == 7'h23 ? _GEN_2282 : DMemory_141; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3307 = EXMEMop == 7'h23 ? _GEN_2283 : DMemory_142; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3308 = EXMEMop == 7'h23 ? _GEN_2284 : DMemory_143; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3309 = EXMEMop == 7'h23 ? _GEN_2285 : DMemory_144; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3310 = EXMEMop == 7'h23 ? _GEN_2286 : DMemory_145; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3311 = EXMEMop == 7'h23 ? _GEN_2287 : DMemory_146; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3312 = EXMEMop == 7'h23 ? _GEN_2288 : DMemory_147; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3313 = EXMEMop == 7'h23 ? _GEN_2289 : DMemory_148; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3314 = EXMEMop == 7'h23 ? _GEN_2290 : DMemory_149; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3315 = EXMEMop == 7'h23 ? _GEN_2291 : DMemory_150; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3316 = EXMEMop == 7'h23 ? _GEN_2292 : DMemory_151; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3317 = EXMEMop == 7'h23 ? _GEN_2293 : DMemory_152; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3318 = EXMEMop == 7'h23 ? _GEN_2294 : DMemory_153; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3319 = EXMEMop == 7'h23 ? _GEN_2295 : DMemory_154; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3320 = EXMEMop == 7'h23 ? _GEN_2296 : DMemory_155; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3321 = EXMEMop == 7'h23 ? _GEN_2297 : DMemory_156; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3322 = EXMEMop == 7'h23 ? _GEN_2298 : DMemory_157; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3323 = EXMEMop == 7'h23 ? _GEN_2299 : DMemory_158; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3324 = EXMEMop == 7'h23 ? _GEN_2300 : DMemory_159; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3325 = EXMEMop == 7'h23 ? _GEN_2301 : DMemory_160; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3326 = EXMEMop == 7'h23 ? _GEN_2302 : DMemory_161; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3327 = EXMEMop == 7'h23 ? _GEN_2303 : DMemory_162; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3328 = EXMEMop == 7'h23 ? _GEN_2304 : DMemory_163; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3329 = EXMEMop == 7'h23 ? _GEN_2305 : DMemory_164; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3330 = EXMEMop == 7'h23 ? _GEN_2306 : DMemory_165; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3331 = EXMEMop == 7'h23 ? _GEN_2307 : DMemory_166; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3332 = EXMEMop == 7'h23 ? _GEN_2308 : DMemory_167; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3333 = EXMEMop == 7'h23 ? _GEN_2309 : DMemory_168; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3334 = EXMEMop == 7'h23 ? _GEN_2310 : DMemory_169; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3335 = EXMEMop == 7'h23 ? _GEN_2311 : DMemory_170; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3336 = EXMEMop == 7'h23 ? _GEN_2312 : DMemory_171; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3337 = EXMEMop == 7'h23 ? _GEN_2313 : DMemory_172; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3338 = EXMEMop == 7'h23 ? _GEN_2314 : DMemory_173; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3339 = EXMEMop == 7'h23 ? _GEN_2315 : DMemory_174; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3340 = EXMEMop == 7'h23 ? _GEN_2316 : DMemory_175; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3341 = EXMEMop == 7'h23 ? _GEN_2317 : DMemory_176; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3342 = EXMEMop == 7'h23 ? _GEN_2318 : DMemory_177; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3343 = EXMEMop == 7'h23 ? _GEN_2319 : DMemory_178; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3344 = EXMEMop == 7'h23 ? _GEN_2320 : DMemory_179; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3345 = EXMEMop == 7'h23 ? _GEN_2321 : DMemory_180; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3346 = EXMEMop == 7'h23 ? _GEN_2322 : DMemory_181; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3347 = EXMEMop == 7'h23 ? _GEN_2323 : DMemory_182; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3348 = EXMEMop == 7'h23 ? _GEN_2324 : DMemory_183; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3349 = EXMEMop == 7'h23 ? _GEN_2325 : DMemory_184; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3350 = EXMEMop == 7'h23 ? _GEN_2326 : DMemory_185; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3351 = EXMEMop == 7'h23 ? _GEN_2327 : DMemory_186; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3352 = EXMEMop == 7'h23 ? _GEN_2328 : DMemory_187; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3353 = EXMEMop == 7'h23 ? _GEN_2329 : DMemory_188; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3354 = EXMEMop == 7'h23 ? _GEN_2330 : DMemory_189; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3355 = EXMEMop == 7'h23 ? _GEN_2331 : DMemory_190; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3356 = EXMEMop == 7'h23 ? _GEN_2332 : DMemory_191; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3357 = EXMEMop == 7'h23 ? _GEN_2333 : DMemory_192; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3358 = EXMEMop == 7'h23 ? _GEN_2334 : DMemory_193; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3359 = EXMEMop == 7'h23 ? _GEN_2335 : DMemory_194; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3360 = EXMEMop == 7'h23 ? _GEN_2336 : DMemory_195; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3361 = EXMEMop == 7'h23 ? _GEN_2337 : DMemory_196; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3362 = EXMEMop == 7'h23 ? _GEN_2338 : DMemory_197; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3363 = EXMEMop == 7'h23 ? _GEN_2339 : DMemory_198; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3364 = EXMEMop == 7'h23 ? _GEN_2340 : DMemory_199; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3365 = EXMEMop == 7'h23 ? _GEN_2341 : DMemory_200; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3366 = EXMEMop == 7'h23 ? _GEN_2342 : DMemory_201; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3367 = EXMEMop == 7'h23 ? _GEN_2343 : DMemory_202; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3368 = EXMEMop == 7'h23 ? _GEN_2344 : DMemory_203; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3369 = EXMEMop == 7'h23 ? _GEN_2345 : DMemory_204; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3370 = EXMEMop == 7'h23 ? _GEN_2346 : DMemory_205; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3371 = EXMEMop == 7'h23 ? _GEN_2347 : DMemory_206; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3372 = EXMEMop == 7'h23 ? _GEN_2348 : DMemory_207; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3373 = EXMEMop == 7'h23 ? _GEN_2349 : DMemory_208; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3374 = EXMEMop == 7'h23 ? _GEN_2350 : DMemory_209; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3375 = EXMEMop == 7'h23 ? _GEN_2351 : DMemory_210; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3376 = EXMEMop == 7'h23 ? _GEN_2352 : DMemory_211; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3377 = EXMEMop == 7'h23 ? _GEN_2353 : DMemory_212; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3378 = EXMEMop == 7'h23 ? _GEN_2354 : DMemory_213; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3379 = EXMEMop == 7'h23 ? _GEN_2355 : DMemory_214; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3380 = EXMEMop == 7'h23 ? _GEN_2356 : DMemory_215; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3381 = EXMEMop == 7'h23 ? _GEN_2357 : DMemory_216; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3382 = EXMEMop == 7'h23 ? _GEN_2358 : DMemory_217; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3383 = EXMEMop == 7'h23 ? _GEN_2359 : DMemory_218; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3384 = EXMEMop == 7'h23 ? _GEN_2360 : DMemory_219; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3385 = EXMEMop == 7'h23 ? _GEN_2361 : DMemory_220; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3386 = EXMEMop == 7'h23 ? _GEN_2362 : DMemory_221; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3387 = EXMEMop == 7'h23 ? _GEN_2363 : DMemory_222; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3388 = EXMEMop == 7'h23 ? _GEN_2364 : DMemory_223; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3389 = EXMEMop == 7'h23 ? _GEN_2365 : DMemory_224; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3390 = EXMEMop == 7'h23 ? _GEN_2366 : DMemory_225; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3391 = EXMEMop == 7'h23 ? _GEN_2367 : DMemory_226; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3392 = EXMEMop == 7'h23 ? _GEN_2368 : DMemory_227; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3393 = EXMEMop == 7'h23 ? _GEN_2369 : DMemory_228; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3394 = EXMEMop == 7'h23 ? _GEN_2370 : DMemory_229; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3395 = EXMEMop == 7'h23 ? _GEN_2371 : DMemory_230; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3396 = EXMEMop == 7'h23 ? _GEN_2372 : DMemory_231; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3397 = EXMEMop == 7'h23 ? _GEN_2373 : DMemory_232; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3398 = EXMEMop == 7'h23 ? _GEN_2374 : DMemory_233; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3399 = EXMEMop == 7'h23 ? _GEN_2375 : DMemory_234; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3400 = EXMEMop == 7'h23 ? _GEN_2376 : DMemory_235; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3401 = EXMEMop == 7'h23 ? _GEN_2377 : DMemory_236; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3402 = EXMEMop == 7'h23 ? _GEN_2378 : DMemory_237; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3403 = EXMEMop == 7'h23 ? _GEN_2379 : DMemory_238; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3404 = EXMEMop == 7'h23 ? _GEN_2380 : DMemory_239; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3405 = EXMEMop == 7'h23 ? _GEN_2381 : DMemory_240; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3406 = EXMEMop == 7'h23 ? _GEN_2382 : DMemory_241; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3407 = EXMEMop == 7'h23 ? _GEN_2383 : DMemory_242; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3408 = EXMEMop == 7'h23 ? _GEN_2384 : DMemory_243; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3409 = EXMEMop == 7'h23 ? _GEN_2385 : DMemory_244; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3410 = EXMEMop == 7'h23 ? _GEN_2386 : DMemory_245; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3411 = EXMEMop == 7'h23 ? _GEN_2387 : DMemory_246; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3412 = EXMEMop == 7'h23 ? _GEN_2388 : DMemory_247; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3413 = EXMEMop == 7'h23 ? _GEN_2389 : DMemory_248; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3414 = EXMEMop == 7'h23 ? _GEN_2390 : DMemory_249; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3415 = EXMEMop == 7'h23 ? _GEN_2391 : DMemory_250; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3416 = EXMEMop == 7'h23 ? _GEN_2392 : DMemory_251; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3417 = EXMEMop == 7'h23 ? _GEN_2393 : DMemory_252; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3418 = EXMEMop == 7'h23 ? _GEN_2394 : DMemory_253; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3419 = EXMEMop == 7'h23 ? _GEN_2395 : DMemory_254; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3420 = EXMEMop == 7'h23 ? _GEN_2396 : DMemory_255; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3421 = EXMEMop == 7'h23 ? _GEN_2397 : DMemory_256; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3422 = EXMEMop == 7'h23 ? _GEN_2398 : DMemory_257; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3423 = EXMEMop == 7'h23 ? _GEN_2399 : DMemory_258; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3424 = EXMEMop == 7'h23 ? _GEN_2400 : DMemory_259; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3425 = EXMEMop == 7'h23 ? _GEN_2401 : DMemory_260; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3426 = EXMEMop == 7'h23 ? _GEN_2402 : DMemory_261; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3427 = EXMEMop == 7'h23 ? _GEN_2403 : DMemory_262; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3428 = EXMEMop == 7'h23 ? _GEN_2404 : DMemory_263; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3429 = EXMEMop == 7'h23 ? _GEN_2405 : DMemory_264; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3430 = EXMEMop == 7'h23 ? _GEN_2406 : DMemory_265; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3431 = EXMEMop == 7'h23 ? _GEN_2407 : DMemory_266; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3432 = EXMEMop == 7'h23 ? _GEN_2408 : DMemory_267; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3433 = EXMEMop == 7'h23 ? _GEN_2409 : DMemory_268; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3434 = EXMEMop == 7'h23 ? _GEN_2410 : DMemory_269; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3435 = EXMEMop == 7'h23 ? _GEN_2411 : DMemory_270; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3436 = EXMEMop == 7'h23 ? _GEN_2412 : DMemory_271; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3437 = EXMEMop == 7'h23 ? _GEN_2413 : DMemory_272; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3438 = EXMEMop == 7'h23 ? _GEN_2414 : DMemory_273; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3439 = EXMEMop == 7'h23 ? _GEN_2415 : DMemory_274; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3440 = EXMEMop == 7'h23 ? _GEN_2416 : DMemory_275; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3441 = EXMEMop == 7'h23 ? _GEN_2417 : DMemory_276; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3442 = EXMEMop == 7'h23 ? _GEN_2418 : DMemory_277; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3443 = EXMEMop == 7'h23 ? _GEN_2419 : DMemory_278; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3444 = EXMEMop == 7'h23 ? _GEN_2420 : DMemory_279; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3445 = EXMEMop == 7'h23 ? _GEN_2421 : DMemory_280; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3446 = EXMEMop == 7'h23 ? _GEN_2422 : DMemory_281; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3447 = EXMEMop == 7'h23 ? _GEN_2423 : DMemory_282; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3448 = EXMEMop == 7'h23 ? _GEN_2424 : DMemory_283; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3449 = EXMEMop == 7'h23 ? _GEN_2425 : DMemory_284; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3450 = EXMEMop == 7'h23 ? _GEN_2426 : DMemory_285; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3451 = EXMEMop == 7'h23 ? _GEN_2427 : DMemory_286; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3452 = EXMEMop == 7'h23 ? _GEN_2428 : DMemory_287; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3453 = EXMEMop == 7'h23 ? _GEN_2429 : DMemory_288; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3454 = EXMEMop == 7'h23 ? _GEN_2430 : DMemory_289; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3455 = EXMEMop == 7'h23 ? _GEN_2431 : DMemory_290; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3456 = EXMEMop == 7'h23 ? _GEN_2432 : DMemory_291; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3457 = EXMEMop == 7'h23 ? _GEN_2433 : DMemory_292; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3458 = EXMEMop == 7'h23 ? _GEN_2434 : DMemory_293; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3459 = EXMEMop == 7'h23 ? _GEN_2435 : DMemory_294; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3460 = EXMEMop == 7'h23 ? _GEN_2436 : DMemory_295; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3461 = EXMEMop == 7'h23 ? _GEN_2437 : DMemory_296; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3462 = EXMEMop == 7'h23 ? _GEN_2438 : DMemory_297; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3463 = EXMEMop == 7'h23 ? _GEN_2439 : DMemory_298; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3464 = EXMEMop == 7'h23 ? _GEN_2440 : DMemory_299; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3465 = EXMEMop == 7'h23 ? _GEN_2441 : DMemory_300; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3466 = EXMEMop == 7'h23 ? _GEN_2442 : DMemory_301; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3467 = EXMEMop == 7'h23 ? _GEN_2443 : DMemory_302; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3468 = EXMEMop == 7'h23 ? _GEN_2444 : DMemory_303; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3469 = EXMEMop == 7'h23 ? _GEN_2445 : DMemory_304; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3470 = EXMEMop == 7'h23 ? _GEN_2446 : DMemory_305; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3471 = EXMEMop == 7'h23 ? _GEN_2447 : DMemory_306; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3472 = EXMEMop == 7'h23 ? _GEN_2448 : DMemory_307; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3473 = EXMEMop == 7'h23 ? _GEN_2449 : DMemory_308; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3474 = EXMEMop == 7'h23 ? _GEN_2450 : DMemory_309; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3475 = EXMEMop == 7'h23 ? _GEN_2451 : DMemory_310; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3476 = EXMEMop == 7'h23 ? _GEN_2452 : DMemory_311; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3477 = EXMEMop == 7'h23 ? _GEN_2453 : DMemory_312; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3478 = EXMEMop == 7'h23 ? _GEN_2454 : DMemory_313; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3479 = EXMEMop == 7'h23 ? _GEN_2455 : DMemory_314; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3480 = EXMEMop == 7'h23 ? _GEN_2456 : DMemory_315; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3481 = EXMEMop == 7'h23 ? _GEN_2457 : DMemory_316; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3482 = EXMEMop == 7'h23 ? _GEN_2458 : DMemory_317; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3483 = EXMEMop == 7'h23 ? _GEN_2459 : DMemory_318; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3484 = EXMEMop == 7'h23 ? _GEN_2460 : DMemory_319; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3485 = EXMEMop == 7'h23 ? _GEN_2461 : DMemory_320; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3486 = EXMEMop == 7'h23 ? _GEN_2462 : DMemory_321; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3487 = EXMEMop == 7'h23 ? _GEN_2463 : DMemory_322; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3488 = EXMEMop == 7'h23 ? _GEN_2464 : DMemory_323; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3489 = EXMEMop == 7'h23 ? _GEN_2465 : DMemory_324; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3490 = EXMEMop == 7'h23 ? _GEN_2466 : DMemory_325; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3491 = EXMEMop == 7'h23 ? _GEN_2467 : DMemory_326; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3492 = EXMEMop == 7'h23 ? _GEN_2468 : DMemory_327; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3493 = EXMEMop == 7'h23 ? _GEN_2469 : DMemory_328; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3494 = EXMEMop == 7'h23 ? _GEN_2470 : DMemory_329; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3495 = EXMEMop == 7'h23 ? _GEN_2471 : DMemory_330; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3496 = EXMEMop == 7'h23 ? _GEN_2472 : DMemory_331; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3497 = EXMEMop == 7'h23 ? _GEN_2473 : DMemory_332; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3498 = EXMEMop == 7'h23 ? _GEN_2474 : DMemory_333; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3499 = EXMEMop == 7'h23 ? _GEN_2475 : DMemory_334; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3500 = EXMEMop == 7'h23 ? _GEN_2476 : DMemory_335; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3501 = EXMEMop == 7'h23 ? _GEN_2477 : DMemory_336; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3502 = EXMEMop == 7'h23 ? _GEN_2478 : DMemory_337; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3503 = EXMEMop == 7'h23 ? _GEN_2479 : DMemory_338; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3504 = EXMEMop == 7'h23 ? _GEN_2480 : DMemory_339; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3505 = EXMEMop == 7'h23 ? _GEN_2481 : DMemory_340; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3506 = EXMEMop == 7'h23 ? _GEN_2482 : DMemory_341; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3507 = EXMEMop == 7'h23 ? _GEN_2483 : DMemory_342; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3508 = EXMEMop == 7'h23 ? _GEN_2484 : DMemory_343; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3509 = EXMEMop == 7'h23 ? _GEN_2485 : DMemory_344; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3510 = EXMEMop == 7'h23 ? _GEN_2486 : DMemory_345; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3511 = EXMEMop == 7'h23 ? _GEN_2487 : DMemory_346; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3512 = EXMEMop == 7'h23 ? _GEN_2488 : DMemory_347; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3513 = EXMEMop == 7'h23 ? _GEN_2489 : DMemory_348; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3514 = EXMEMop == 7'h23 ? _GEN_2490 : DMemory_349; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3515 = EXMEMop == 7'h23 ? _GEN_2491 : DMemory_350; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3516 = EXMEMop == 7'h23 ? _GEN_2492 : DMemory_351; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3517 = EXMEMop == 7'h23 ? _GEN_2493 : DMemory_352; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3518 = EXMEMop == 7'h23 ? _GEN_2494 : DMemory_353; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3519 = EXMEMop == 7'h23 ? _GEN_2495 : DMemory_354; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3520 = EXMEMop == 7'h23 ? _GEN_2496 : DMemory_355; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3521 = EXMEMop == 7'h23 ? _GEN_2497 : DMemory_356; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3522 = EXMEMop == 7'h23 ? _GEN_2498 : DMemory_357; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3523 = EXMEMop == 7'h23 ? _GEN_2499 : DMemory_358; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3524 = EXMEMop == 7'h23 ? _GEN_2500 : DMemory_359; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3525 = EXMEMop == 7'h23 ? _GEN_2501 : DMemory_360; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3526 = EXMEMop == 7'h23 ? _GEN_2502 : DMemory_361; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3527 = EXMEMop == 7'h23 ? _GEN_2503 : DMemory_362; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3528 = EXMEMop == 7'h23 ? _GEN_2504 : DMemory_363; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3529 = EXMEMop == 7'h23 ? _GEN_2505 : DMemory_364; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3530 = EXMEMop == 7'h23 ? _GEN_2506 : DMemory_365; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3531 = EXMEMop == 7'h23 ? _GEN_2507 : DMemory_366; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3532 = EXMEMop == 7'h23 ? _GEN_2508 : DMemory_367; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3533 = EXMEMop == 7'h23 ? _GEN_2509 : DMemory_368; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3534 = EXMEMop == 7'h23 ? _GEN_2510 : DMemory_369; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3535 = EXMEMop == 7'h23 ? _GEN_2511 : DMemory_370; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3536 = EXMEMop == 7'h23 ? _GEN_2512 : DMemory_371; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3537 = EXMEMop == 7'h23 ? _GEN_2513 : DMemory_372; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3538 = EXMEMop == 7'h23 ? _GEN_2514 : DMemory_373; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3539 = EXMEMop == 7'h23 ? _GEN_2515 : DMemory_374; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3540 = EXMEMop == 7'h23 ? _GEN_2516 : DMemory_375; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3541 = EXMEMop == 7'h23 ? _GEN_2517 : DMemory_376; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3542 = EXMEMop == 7'h23 ? _GEN_2518 : DMemory_377; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3543 = EXMEMop == 7'h23 ? _GEN_2519 : DMemory_378; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3544 = EXMEMop == 7'h23 ? _GEN_2520 : DMemory_379; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3545 = EXMEMop == 7'h23 ? _GEN_2521 : DMemory_380; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3546 = EXMEMop == 7'h23 ? _GEN_2522 : DMemory_381; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3547 = EXMEMop == 7'h23 ? _GEN_2523 : DMemory_382; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3548 = EXMEMop == 7'h23 ? _GEN_2524 : DMemory_383; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3549 = EXMEMop == 7'h23 ? _GEN_2525 : DMemory_384; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3550 = EXMEMop == 7'h23 ? _GEN_2526 : DMemory_385; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3551 = EXMEMop == 7'h23 ? _GEN_2527 : DMemory_386; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3552 = EXMEMop == 7'h23 ? _GEN_2528 : DMemory_387; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3553 = EXMEMop == 7'h23 ? _GEN_2529 : DMemory_388; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3554 = EXMEMop == 7'h23 ? _GEN_2530 : DMemory_389; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3555 = EXMEMop == 7'h23 ? _GEN_2531 : DMemory_390; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3556 = EXMEMop == 7'h23 ? _GEN_2532 : DMemory_391; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3557 = EXMEMop == 7'h23 ? _GEN_2533 : DMemory_392; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3558 = EXMEMop == 7'h23 ? _GEN_2534 : DMemory_393; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3559 = EXMEMop == 7'h23 ? _GEN_2535 : DMemory_394; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3560 = EXMEMop == 7'h23 ? _GEN_2536 : DMemory_395; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3561 = EXMEMop == 7'h23 ? _GEN_2537 : DMemory_396; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3562 = EXMEMop == 7'h23 ? _GEN_2538 : DMemory_397; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3563 = EXMEMop == 7'h23 ? _GEN_2539 : DMemory_398; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3564 = EXMEMop == 7'h23 ? _GEN_2540 : DMemory_399; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3565 = EXMEMop == 7'h23 ? _GEN_2541 : DMemory_400; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3566 = EXMEMop == 7'h23 ? _GEN_2542 : DMemory_401; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3567 = EXMEMop == 7'h23 ? _GEN_2543 : DMemory_402; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3568 = EXMEMop == 7'h23 ? _GEN_2544 : DMemory_403; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3569 = EXMEMop == 7'h23 ? _GEN_2545 : DMemory_404; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3570 = EXMEMop == 7'h23 ? _GEN_2546 : DMemory_405; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3571 = EXMEMop == 7'h23 ? _GEN_2547 : DMemory_406; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3572 = EXMEMop == 7'h23 ? _GEN_2548 : DMemory_407; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3573 = EXMEMop == 7'h23 ? _GEN_2549 : DMemory_408; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3574 = EXMEMop == 7'h23 ? _GEN_2550 : DMemory_409; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3575 = EXMEMop == 7'h23 ? _GEN_2551 : DMemory_410; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3576 = EXMEMop == 7'h23 ? _GEN_2552 : DMemory_411; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3577 = EXMEMop == 7'h23 ? _GEN_2553 : DMemory_412; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3578 = EXMEMop == 7'h23 ? _GEN_2554 : DMemory_413; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3579 = EXMEMop == 7'h23 ? _GEN_2555 : DMemory_414; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3580 = EXMEMop == 7'h23 ? _GEN_2556 : DMemory_415; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3581 = EXMEMop == 7'h23 ? _GEN_2557 : DMemory_416; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3582 = EXMEMop == 7'h23 ? _GEN_2558 : DMemory_417; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3583 = EXMEMop == 7'h23 ? _GEN_2559 : DMemory_418; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3584 = EXMEMop == 7'h23 ? _GEN_2560 : DMemory_419; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3585 = EXMEMop == 7'h23 ? _GEN_2561 : DMemory_420; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3586 = EXMEMop == 7'h23 ? _GEN_2562 : DMemory_421; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3587 = EXMEMop == 7'h23 ? _GEN_2563 : DMemory_422; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3588 = EXMEMop == 7'h23 ? _GEN_2564 : DMemory_423; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3589 = EXMEMop == 7'h23 ? _GEN_2565 : DMemory_424; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3590 = EXMEMop == 7'h23 ? _GEN_2566 : DMemory_425; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3591 = EXMEMop == 7'h23 ? _GEN_2567 : DMemory_426; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3592 = EXMEMop == 7'h23 ? _GEN_2568 : DMemory_427; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3593 = EXMEMop == 7'h23 ? _GEN_2569 : DMemory_428; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3594 = EXMEMop == 7'h23 ? _GEN_2570 : DMemory_429; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3595 = EXMEMop == 7'h23 ? _GEN_2571 : DMemory_430; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3596 = EXMEMop == 7'h23 ? _GEN_2572 : DMemory_431; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3597 = EXMEMop == 7'h23 ? _GEN_2573 : DMemory_432; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3598 = EXMEMop == 7'h23 ? _GEN_2574 : DMemory_433; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3599 = EXMEMop == 7'h23 ? _GEN_2575 : DMemory_434; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3600 = EXMEMop == 7'h23 ? _GEN_2576 : DMemory_435; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3601 = EXMEMop == 7'h23 ? _GEN_2577 : DMemory_436; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3602 = EXMEMop == 7'h23 ? _GEN_2578 : DMemory_437; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3603 = EXMEMop == 7'h23 ? _GEN_2579 : DMemory_438; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3604 = EXMEMop == 7'h23 ? _GEN_2580 : DMemory_439; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3605 = EXMEMop == 7'h23 ? _GEN_2581 : DMemory_440; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3606 = EXMEMop == 7'h23 ? _GEN_2582 : DMemory_441; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3607 = EXMEMop == 7'h23 ? _GEN_2583 : DMemory_442; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3608 = EXMEMop == 7'h23 ? _GEN_2584 : DMemory_443; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3609 = EXMEMop == 7'h23 ? _GEN_2585 : DMemory_444; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3610 = EXMEMop == 7'h23 ? _GEN_2586 : DMemory_445; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3611 = EXMEMop == 7'h23 ? _GEN_2587 : DMemory_446; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3612 = EXMEMop == 7'h23 ? _GEN_2588 : DMemory_447; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3613 = EXMEMop == 7'h23 ? _GEN_2589 : DMemory_448; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3614 = EXMEMop == 7'h23 ? _GEN_2590 : DMemory_449; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3615 = EXMEMop == 7'h23 ? _GEN_2591 : DMemory_450; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3616 = EXMEMop == 7'h23 ? _GEN_2592 : DMemory_451; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3617 = EXMEMop == 7'h23 ? _GEN_2593 : DMemory_452; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3618 = EXMEMop == 7'h23 ? _GEN_2594 : DMemory_453; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3619 = EXMEMop == 7'h23 ? _GEN_2595 : DMemory_454; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3620 = EXMEMop == 7'h23 ? _GEN_2596 : DMemory_455; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3621 = EXMEMop == 7'h23 ? _GEN_2597 : DMemory_456; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3622 = EXMEMop == 7'h23 ? _GEN_2598 : DMemory_457; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3623 = EXMEMop == 7'h23 ? _GEN_2599 : DMemory_458; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3624 = EXMEMop == 7'h23 ? _GEN_2600 : DMemory_459; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3625 = EXMEMop == 7'h23 ? _GEN_2601 : DMemory_460; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3626 = EXMEMop == 7'h23 ? _GEN_2602 : DMemory_461; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3627 = EXMEMop == 7'h23 ? _GEN_2603 : DMemory_462; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3628 = EXMEMop == 7'h23 ? _GEN_2604 : DMemory_463; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3629 = EXMEMop == 7'h23 ? _GEN_2605 : DMemory_464; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3630 = EXMEMop == 7'h23 ? _GEN_2606 : DMemory_465; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3631 = EXMEMop == 7'h23 ? _GEN_2607 : DMemory_466; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3632 = EXMEMop == 7'h23 ? _GEN_2608 : DMemory_467; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3633 = EXMEMop == 7'h23 ? _GEN_2609 : DMemory_468; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3634 = EXMEMop == 7'h23 ? _GEN_2610 : DMemory_469; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3635 = EXMEMop == 7'h23 ? _GEN_2611 : DMemory_470; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3636 = EXMEMop == 7'h23 ? _GEN_2612 : DMemory_471; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3637 = EXMEMop == 7'h23 ? _GEN_2613 : DMemory_472; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3638 = EXMEMop == 7'h23 ? _GEN_2614 : DMemory_473; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3639 = EXMEMop == 7'h23 ? _GEN_2615 : DMemory_474; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3640 = EXMEMop == 7'h23 ? _GEN_2616 : DMemory_475; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3641 = EXMEMop == 7'h23 ? _GEN_2617 : DMemory_476; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3642 = EXMEMop == 7'h23 ? _GEN_2618 : DMemory_477; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3643 = EXMEMop == 7'h23 ? _GEN_2619 : DMemory_478; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3644 = EXMEMop == 7'h23 ? _GEN_2620 : DMemory_479; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3645 = EXMEMop == 7'h23 ? _GEN_2621 : DMemory_480; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3646 = EXMEMop == 7'h23 ? _GEN_2622 : DMemory_481; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3647 = EXMEMop == 7'h23 ? _GEN_2623 : DMemory_482; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3648 = EXMEMop == 7'h23 ? _GEN_2624 : DMemory_483; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3649 = EXMEMop == 7'h23 ? _GEN_2625 : DMemory_484; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3650 = EXMEMop == 7'h23 ? _GEN_2626 : DMemory_485; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3651 = EXMEMop == 7'h23 ? _GEN_2627 : DMemory_486; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3652 = EXMEMop == 7'h23 ? _GEN_2628 : DMemory_487; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3653 = EXMEMop == 7'h23 ? _GEN_2629 : DMemory_488; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3654 = EXMEMop == 7'h23 ? _GEN_2630 : DMemory_489; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3655 = EXMEMop == 7'h23 ? _GEN_2631 : DMemory_490; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3656 = EXMEMop == 7'h23 ? _GEN_2632 : DMemory_491; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3657 = EXMEMop == 7'h23 ? _GEN_2633 : DMemory_492; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3658 = EXMEMop == 7'h23 ? _GEN_2634 : DMemory_493; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3659 = EXMEMop == 7'h23 ? _GEN_2635 : DMemory_494; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3660 = EXMEMop == 7'h23 ? _GEN_2636 : DMemory_495; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3661 = EXMEMop == 7'h23 ? _GEN_2637 : DMemory_496; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3662 = EXMEMop == 7'h23 ? _GEN_2638 : DMemory_497; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3663 = EXMEMop == 7'h23 ? _GEN_2639 : DMemory_498; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3664 = EXMEMop == 7'h23 ? _GEN_2640 : DMemory_499; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3665 = EXMEMop == 7'h23 ? _GEN_2641 : DMemory_500; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3666 = EXMEMop == 7'h23 ? _GEN_2642 : DMemory_501; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3667 = EXMEMop == 7'h23 ? _GEN_2643 : DMemory_502; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3668 = EXMEMop == 7'h23 ? _GEN_2644 : DMemory_503; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3669 = EXMEMop == 7'h23 ? _GEN_2645 : DMemory_504; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3670 = EXMEMop == 7'h23 ? _GEN_2646 : DMemory_505; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3671 = EXMEMop == 7'h23 ? _GEN_2647 : DMemory_506; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3672 = EXMEMop == 7'h23 ? _GEN_2648 : DMemory_507; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3673 = EXMEMop == 7'h23 ? _GEN_2649 : DMemory_508; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3674 = EXMEMop == 7'h23 ? _GEN_2650 : DMemory_509; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3675 = EXMEMop == 7'h23 ? _GEN_2651 : DMemory_510; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3676 = EXMEMop == 7'h23 ? _GEN_2652 : DMemory_511; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3677 = EXMEMop == 7'h23 ? _GEN_2653 : DMemory_512; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3678 = EXMEMop == 7'h23 ? _GEN_2654 : DMemory_513; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3679 = EXMEMop == 7'h23 ? _GEN_2655 : DMemory_514; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3680 = EXMEMop == 7'h23 ? _GEN_2656 : DMemory_515; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3681 = EXMEMop == 7'h23 ? _GEN_2657 : DMemory_516; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3682 = EXMEMop == 7'h23 ? _GEN_2658 : DMemory_517; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3683 = EXMEMop == 7'h23 ? _GEN_2659 : DMemory_518; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3684 = EXMEMop == 7'h23 ? _GEN_2660 : DMemory_519; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3685 = EXMEMop == 7'h23 ? _GEN_2661 : DMemory_520; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3686 = EXMEMop == 7'h23 ? _GEN_2662 : DMemory_521; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3687 = EXMEMop == 7'h23 ? _GEN_2663 : DMemory_522; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3688 = EXMEMop == 7'h23 ? _GEN_2664 : DMemory_523; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3689 = EXMEMop == 7'h23 ? _GEN_2665 : DMemory_524; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3690 = EXMEMop == 7'h23 ? _GEN_2666 : DMemory_525; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3691 = EXMEMop == 7'h23 ? _GEN_2667 : DMemory_526; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3692 = EXMEMop == 7'h23 ? _GEN_2668 : DMemory_527; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3693 = EXMEMop == 7'h23 ? _GEN_2669 : DMemory_528; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3694 = EXMEMop == 7'h23 ? _GEN_2670 : DMemory_529; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3695 = EXMEMop == 7'h23 ? _GEN_2671 : DMemory_530; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3696 = EXMEMop == 7'h23 ? _GEN_2672 : DMemory_531; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3697 = EXMEMop == 7'h23 ? _GEN_2673 : DMemory_532; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3698 = EXMEMop == 7'h23 ? _GEN_2674 : DMemory_533; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3699 = EXMEMop == 7'h23 ? _GEN_2675 : DMemory_534; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3700 = EXMEMop == 7'h23 ? _GEN_2676 : DMemory_535; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3701 = EXMEMop == 7'h23 ? _GEN_2677 : DMemory_536; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3702 = EXMEMop == 7'h23 ? _GEN_2678 : DMemory_537; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3703 = EXMEMop == 7'h23 ? _GEN_2679 : DMemory_538; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3704 = EXMEMop == 7'h23 ? _GEN_2680 : DMemory_539; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3705 = EXMEMop == 7'h23 ? _GEN_2681 : DMemory_540; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3706 = EXMEMop == 7'h23 ? _GEN_2682 : DMemory_541; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3707 = EXMEMop == 7'h23 ? _GEN_2683 : DMemory_542; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3708 = EXMEMop == 7'h23 ? _GEN_2684 : DMemory_543; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3709 = EXMEMop == 7'h23 ? _GEN_2685 : DMemory_544; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3710 = EXMEMop == 7'h23 ? _GEN_2686 : DMemory_545; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3711 = EXMEMop == 7'h23 ? _GEN_2687 : DMemory_546; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3712 = EXMEMop == 7'h23 ? _GEN_2688 : DMemory_547; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3713 = EXMEMop == 7'h23 ? _GEN_2689 : DMemory_548; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3714 = EXMEMop == 7'h23 ? _GEN_2690 : DMemory_549; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3715 = EXMEMop == 7'h23 ? _GEN_2691 : DMemory_550; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3716 = EXMEMop == 7'h23 ? _GEN_2692 : DMemory_551; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3717 = EXMEMop == 7'h23 ? _GEN_2693 : DMemory_552; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3718 = EXMEMop == 7'h23 ? _GEN_2694 : DMemory_553; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3719 = EXMEMop == 7'h23 ? _GEN_2695 : DMemory_554; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3720 = EXMEMop == 7'h23 ? _GEN_2696 : DMemory_555; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3721 = EXMEMop == 7'h23 ? _GEN_2697 : DMemory_556; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3722 = EXMEMop == 7'h23 ? _GEN_2698 : DMemory_557; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3723 = EXMEMop == 7'h23 ? _GEN_2699 : DMemory_558; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3724 = EXMEMop == 7'h23 ? _GEN_2700 : DMemory_559; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3725 = EXMEMop == 7'h23 ? _GEN_2701 : DMemory_560; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3726 = EXMEMop == 7'h23 ? _GEN_2702 : DMemory_561; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3727 = EXMEMop == 7'h23 ? _GEN_2703 : DMemory_562; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3728 = EXMEMop == 7'h23 ? _GEN_2704 : DMemory_563; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3729 = EXMEMop == 7'h23 ? _GEN_2705 : DMemory_564; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3730 = EXMEMop == 7'h23 ? _GEN_2706 : DMemory_565; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3731 = EXMEMop == 7'h23 ? _GEN_2707 : DMemory_566; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3732 = EXMEMop == 7'h23 ? _GEN_2708 : DMemory_567; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3733 = EXMEMop == 7'h23 ? _GEN_2709 : DMemory_568; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3734 = EXMEMop == 7'h23 ? _GEN_2710 : DMemory_569; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3735 = EXMEMop == 7'h23 ? _GEN_2711 : DMemory_570; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3736 = EXMEMop == 7'h23 ? _GEN_2712 : DMemory_571; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3737 = EXMEMop == 7'h23 ? _GEN_2713 : DMemory_572; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3738 = EXMEMop == 7'h23 ? _GEN_2714 : DMemory_573; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3739 = EXMEMop == 7'h23 ? _GEN_2715 : DMemory_574; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3740 = EXMEMop == 7'h23 ? _GEN_2716 : DMemory_575; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3741 = EXMEMop == 7'h23 ? _GEN_2717 : DMemory_576; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3742 = EXMEMop == 7'h23 ? _GEN_2718 : DMemory_577; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3743 = EXMEMop == 7'h23 ? _GEN_2719 : DMemory_578; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3744 = EXMEMop == 7'h23 ? _GEN_2720 : DMemory_579; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3745 = EXMEMop == 7'h23 ? _GEN_2721 : DMemory_580; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3746 = EXMEMop == 7'h23 ? _GEN_2722 : DMemory_581; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3747 = EXMEMop == 7'h23 ? _GEN_2723 : DMemory_582; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3748 = EXMEMop == 7'h23 ? _GEN_2724 : DMemory_583; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3749 = EXMEMop == 7'h23 ? _GEN_2725 : DMemory_584; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3750 = EXMEMop == 7'h23 ? _GEN_2726 : DMemory_585; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3751 = EXMEMop == 7'h23 ? _GEN_2727 : DMemory_586; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3752 = EXMEMop == 7'h23 ? _GEN_2728 : DMemory_587; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3753 = EXMEMop == 7'h23 ? _GEN_2729 : DMemory_588; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3754 = EXMEMop == 7'h23 ? _GEN_2730 : DMemory_589; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3755 = EXMEMop == 7'h23 ? _GEN_2731 : DMemory_590; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3756 = EXMEMop == 7'h23 ? _GEN_2732 : DMemory_591; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3757 = EXMEMop == 7'h23 ? _GEN_2733 : DMemory_592; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3758 = EXMEMop == 7'h23 ? _GEN_2734 : DMemory_593; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3759 = EXMEMop == 7'h23 ? _GEN_2735 : DMemory_594; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3760 = EXMEMop == 7'h23 ? _GEN_2736 : DMemory_595; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3761 = EXMEMop == 7'h23 ? _GEN_2737 : DMemory_596; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3762 = EXMEMop == 7'h23 ? _GEN_2738 : DMemory_597; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3763 = EXMEMop == 7'h23 ? _GEN_2739 : DMemory_598; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3764 = EXMEMop == 7'h23 ? _GEN_2740 : DMemory_599; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3765 = EXMEMop == 7'h23 ? _GEN_2741 : DMemory_600; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3766 = EXMEMop == 7'h23 ? _GEN_2742 : DMemory_601; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3767 = EXMEMop == 7'h23 ? _GEN_2743 : DMemory_602; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3768 = EXMEMop == 7'h23 ? _GEN_2744 : DMemory_603; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3769 = EXMEMop == 7'h23 ? _GEN_2745 : DMemory_604; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3770 = EXMEMop == 7'h23 ? _GEN_2746 : DMemory_605; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3771 = EXMEMop == 7'h23 ? _GEN_2747 : DMemory_606; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3772 = EXMEMop == 7'h23 ? _GEN_2748 : DMemory_607; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3773 = EXMEMop == 7'h23 ? _GEN_2749 : DMemory_608; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3774 = EXMEMop == 7'h23 ? _GEN_2750 : DMemory_609; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3775 = EXMEMop == 7'h23 ? _GEN_2751 : DMemory_610; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3776 = EXMEMop == 7'h23 ? _GEN_2752 : DMemory_611; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3777 = EXMEMop == 7'h23 ? _GEN_2753 : DMemory_612; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3778 = EXMEMop == 7'h23 ? _GEN_2754 : DMemory_613; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3779 = EXMEMop == 7'h23 ? _GEN_2755 : DMemory_614; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3780 = EXMEMop == 7'h23 ? _GEN_2756 : DMemory_615; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3781 = EXMEMop == 7'h23 ? _GEN_2757 : DMemory_616; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3782 = EXMEMop == 7'h23 ? _GEN_2758 : DMemory_617; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3783 = EXMEMop == 7'h23 ? _GEN_2759 : DMemory_618; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3784 = EXMEMop == 7'h23 ? _GEN_2760 : DMemory_619; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3785 = EXMEMop == 7'h23 ? _GEN_2761 : DMemory_620; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3786 = EXMEMop == 7'h23 ? _GEN_2762 : DMemory_621; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3787 = EXMEMop == 7'h23 ? _GEN_2763 : DMemory_622; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3788 = EXMEMop == 7'h23 ? _GEN_2764 : DMemory_623; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3789 = EXMEMop == 7'h23 ? _GEN_2765 : DMemory_624; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3790 = EXMEMop == 7'h23 ? _GEN_2766 : DMemory_625; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3791 = EXMEMop == 7'h23 ? _GEN_2767 : DMemory_626; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3792 = EXMEMop == 7'h23 ? _GEN_2768 : DMemory_627; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3793 = EXMEMop == 7'h23 ? _GEN_2769 : DMemory_628; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3794 = EXMEMop == 7'h23 ? _GEN_2770 : DMemory_629; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3795 = EXMEMop == 7'h23 ? _GEN_2771 : DMemory_630; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3796 = EXMEMop == 7'h23 ? _GEN_2772 : DMemory_631; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3797 = EXMEMop == 7'h23 ? _GEN_2773 : DMemory_632; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3798 = EXMEMop == 7'h23 ? _GEN_2774 : DMemory_633; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3799 = EXMEMop == 7'h23 ? _GEN_2775 : DMemory_634; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3800 = EXMEMop == 7'h23 ? _GEN_2776 : DMemory_635; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3801 = EXMEMop == 7'h23 ? _GEN_2777 : DMemory_636; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3802 = EXMEMop == 7'h23 ? _GEN_2778 : DMemory_637; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3803 = EXMEMop == 7'h23 ? _GEN_2779 : DMemory_638; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3804 = EXMEMop == 7'h23 ? _GEN_2780 : DMemory_639; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3805 = EXMEMop == 7'h23 ? _GEN_2781 : DMemory_640; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3806 = EXMEMop == 7'h23 ? _GEN_2782 : DMemory_641; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3807 = EXMEMop == 7'h23 ? _GEN_2783 : DMemory_642; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3808 = EXMEMop == 7'h23 ? _GEN_2784 : DMemory_643; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3809 = EXMEMop == 7'h23 ? _GEN_2785 : DMemory_644; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3810 = EXMEMop == 7'h23 ? _GEN_2786 : DMemory_645; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3811 = EXMEMop == 7'h23 ? _GEN_2787 : DMemory_646; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3812 = EXMEMop == 7'h23 ? _GEN_2788 : DMemory_647; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3813 = EXMEMop == 7'h23 ? _GEN_2789 : DMemory_648; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3814 = EXMEMop == 7'h23 ? _GEN_2790 : DMemory_649; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3815 = EXMEMop == 7'h23 ? _GEN_2791 : DMemory_650; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3816 = EXMEMop == 7'h23 ? _GEN_2792 : DMemory_651; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3817 = EXMEMop == 7'h23 ? _GEN_2793 : DMemory_652; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3818 = EXMEMop == 7'h23 ? _GEN_2794 : DMemory_653; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3819 = EXMEMop == 7'h23 ? _GEN_2795 : DMemory_654; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3820 = EXMEMop == 7'h23 ? _GEN_2796 : DMemory_655; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3821 = EXMEMop == 7'h23 ? _GEN_2797 : DMemory_656; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3822 = EXMEMop == 7'h23 ? _GEN_2798 : DMemory_657; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3823 = EXMEMop == 7'h23 ? _GEN_2799 : DMemory_658; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3824 = EXMEMop == 7'h23 ? _GEN_2800 : DMemory_659; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3825 = EXMEMop == 7'h23 ? _GEN_2801 : DMemory_660; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3826 = EXMEMop == 7'h23 ? _GEN_2802 : DMemory_661; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3827 = EXMEMop == 7'h23 ? _GEN_2803 : DMemory_662; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3828 = EXMEMop == 7'h23 ? _GEN_2804 : DMemory_663; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3829 = EXMEMop == 7'h23 ? _GEN_2805 : DMemory_664; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3830 = EXMEMop == 7'h23 ? _GEN_2806 : DMemory_665; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3831 = EXMEMop == 7'h23 ? _GEN_2807 : DMemory_666; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3832 = EXMEMop == 7'h23 ? _GEN_2808 : DMemory_667; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3833 = EXMEMop == 7'h23 ? _GEN_2809 : DMemory_668; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3834 = EXMEMop == 7'h23 ? _GEN_2810 : DMemory_669; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3835 = EXMEMop == 7'h23 ? _GEN_2811 : DMemory_670; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3836 = EXMEMop == 7'h23 ? _GEN_2812 : DMemory_671; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3837 = EXMEMop == 7'h23 ? _GEN_2813 : DMemory_672; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3838 = EXMEMop == 7'h23 ? _GEN_2814 : DMemory_673; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3839 = EXMEMop == 7'h23 ? _GEN_2815 : DMemory_674; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3840 = EXMEMop == 7'h23 ? _GEN_2816 : DMemory_675; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3841 = EXMEMop == 7'h23 ? _GEN_2817 : DMemory_676; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3842 = EXMEMop == 7'h23 ? _GEN_2818 : DMemory_677; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3843 = EXMEMop == 7'h23 ? _GEN_2819 : DMemory_678; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3844 = EXMEMop == 7'h23 ? _GEN_2820 : DMemory_679; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3845 = EXMEMop == 7'h23 ? _GEN_2821 : DMemory_680; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3846 = EXMEMop == 7'h23 ? _GEN_2822 : DMemory_681; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3847 = EXMEMop == 7'h23 ? _GEN_2823 : DMemory_682; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3848 = EXMEMop == 7'h23 ? _GEN_2824 : DMemory_683; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3849 = EXMEMop == 7'h23 ? _GEN_2825 : DMemory_684; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3850 = EXMEMop == 7'h23 ? _GEN_2826 : DMemory_685; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3851 = EXMEMop == 7'h23 ? _GEN_2827 : DMemory_686; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3852 = EXMEMop == 7'h23 ? _GEN_2828 : DMemory_687; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3853 = EXMEMop == 7'h23 ? _GEN_2829 : DMemory_688; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3854 = EXMEMop == 7'h23 ? _GEN_2830 : DMemory_689; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3855 = EXMEMop == 7'h23 ? _GEN_2831 : DMemory_690; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3856 = EXMEMop == 7'h23 ? _GEN_2832 : DMemory_691; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3857 = EXMEMop == 7'h23 ? _GEN_2833 : DMemory_692; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3858 = EXMEMop == 7'h23 ? _GEN_2834 : DMemory_693; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3859 = EXMEMop == 7'h23 ? _GEN_2835 : DMemory_694; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3860 = EXMEMop == 7'h23 ? _GEN_2836 : DMemory_695; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3861 = EXMEMop == 7'h23 ? _GEN_2837 : DMemory_696; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3862 = EXMEMop == 7'h23 ? _GEN_2838 : DMemory_697; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3863 = EXMEMop == 7'h23 ? _GEN_2839 : DMemory_698; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3864 = EXMEMop == 7'h23 ? _GEN_2840 : DMemory_699; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3865 = EXMEMop == 7'h23 ? _GEN_2841 : DMemory_700; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3866 = EXMEMop == 7'h23 ? _GEN_2842 : DMemory_701; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3867 = EXMEMop == 7'h23 ? _GEN_2843 : DMemory_702; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3868 = EXMEMop == 7'h23 ? _GEN_2844 : DMemory_703; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3869 = EXMEMop == 7'h23 ? _GEN_2845 : DMemory_704; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3870 = EXMEMop == 7'h23 ? _GEN_2846 : DMemory_705; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3871 = EXMEMop == 7'h23 ? _GEN_2847 : DMemory_706; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3872 = EXMEMop == 7'h23 ? _GEN_2848 : DMemory_707; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3873 = EXMEMop == 7'h23 ? _GEN_2849 : DMemory_708; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3874 = EXMEMop == 7'h23 ? _GEN_2850 : DMemory_709; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3875 = EXMEMop == 7'h23 ? _GEN_2851 : DMemory_710; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3876 = EXMEMop == 7'h23 ? _GEN_2852 : DMemory_711; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3877 = EXMEMop == 7'h23 ? _GEN_2853 : DMemory_712; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3878 = EXMEMop == 7'h23 ? _GEN_2854 : DMemory_713; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3879 = EXMEMop == 7'h23 ? _GEN_2855 : DMemory_714; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3880 = EXMEMop == 7'h23 ? _GEN_2856 : DMemory_715; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3881 = EXMEMop == 7'h23 ? _GEN_2857 : DMemory_716; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3882 = EXMEMop == 7'h23 ? _GEN_2858 : DMemory_717; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3883 = EXMEMop == 7'h23 ? _GEN_2859 : DMemory_718; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3884 = EXMEMop == 7'h23 ? _GEN_2860 : DMemory_719; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3885 = EXMEMop == 7'h23 ? _GEN_2861 : DMemory_720; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3886 = EXMEMop == 7'h23 ? _GEN_2862 : DMemory_721; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3887 = EXMEMop == 7'h23 ? _GEN_2863 : DMemory_722; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3888 = EXMEMop == 7'h23 ? _GEN_2864 : DMemory_723; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3889 = EXMEMop == 7'h23 ? _GEN_2865 : DMemory_724; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3890 = EXMEMop == 7'h23 ? _GEN_2866 : DMemory_725; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3891 = EXMEMop == 7'h23 ? _GEN_2867 : DMemory_726; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3892 = EXMEMop == 7'h23 ? _GEN_2868 : DMemory_727; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3893 = EXMEMop == 7'h23 ? _GEN_2869 : DMemory_728; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3894 = EXMEMop == 7'h23 ? _GEN_2870 : DMemory_729; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3895 = EXMEMop == 7'h23 ? _GEN_2871 : DMemory_730; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3896 = EXMEMop == 7'h23 ? _GEN_2872 : DMemory_731; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3897 = EXMEMop == 7'h23 ? _GEN_2873 : DMemory_732; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3898 = EXMEMop == 7'h23 ? _GEN_2874 : DMemory_733; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3899 = EXMEMop == 7'h23 ? _GEN_2875 : DMemory_734; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3900 = EXMEMop == 7'h23 ? _GEN_2876 : DMemory_735; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3901 = EXMEMop == 7'h23 ? _GEN_2877 : DMemory_736; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3902 = EXMEMop == 7'h23 ? _GEN_2878 : DMemory_737; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3903 = EXMEMop == 7'h23 ? _GEN_2879 : DMemory_738; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3904 = EXMEMop == 7'h23 ? _GEN_2880 : DMemory_739; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3905 = EXMEMop == 7'h23 ? _GEN_2881 : DMemory_740; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3906 = EXMEMop == 7'h23 ? _GEN_2882 : DMemory_741; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3907 = EXMEMop == 7'h23 ? _GEN_2883 : DMemory_742; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3908 = EXMEMop == 7'h23 ? _GEN_2884 : DMemory_743; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3909 = EXMEMop == 7'h23 ? _GEN_2885 : DMemory_744; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3910 = EXMEMop == 7'h23 ? _GEN_2886 : DMemory_745; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3911 = EXMEMop == 7'h23 ? _GEN_2887 : DMemory_746; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3912 = EXMEMop == 7'h23 ? _GEN_2888 : DMemory_747; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3913 = EXMEMop == 7'h23 ? _GEN_2889 : DMemory_748; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3914 = EXMEMop == 7'h23 ? _GEN_2890 : DMemory_749; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3915 = EXMEMop == 7'h23 ? _GEN_2891 : DMemory_750; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3916 = EXMEMop == 7'h23 ? _GEN_2892 : DMemory_751; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3917 = EXMEMop == 7'h23 ? _GEN_2893 : DMemory_752; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3918 = EXMEMop == 7'h23 ? _GEN_2894 : DMemory_753; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3919 = EXMEMop == 7'h23 ? _GEN_2895 : DMemory_754; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3920 = EXMEMop == 7'h23 ? _GEN_2896 : DMemory_755; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3921 = EXMEMop == 7'h23 ? _GEN_2897 : DMemory_756; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3922 = EXMEMop == 7'h23 ? _GEN_2898 : DMemory_757; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3923 = EXMEMop == 7'h23 ? _GEN_2899 : DMemory_758; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3924 = EXMEMop == 7'h23 ? _GEN_2900 : DMemory_759; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3925 = EXMEMop == 7'h23 ? _GEN_2901 : DMemory_760; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3926 = EXMEMop == 7'h23 ? _GEN_2902 : DMemory_761; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3927 = EXMEMop == 7'h23 ? _GEN_2903 : DMemory_762; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3928 = EXMEMop == 7'h23 ? _GEN_2904 : DMemory_763; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3929 = EXMEMop == 7'h23 ? _GEN_2905 : DMemory_764; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3930 = EXMEMop == 7'h23 ? _GEN_2906 : DMemory_765; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3931 = EXMEMop == 7'h23 ? _GEN_2907 : DMemory_766; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3932 = EXMEMop == 7'h23 ? _GEN_2908 : DMemory_767; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3933 = EXMEMop == 7'h23 ? _GEN_2909 : DMemory_768; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3934 = EXMEMop == 7'h23 ? _GEN_2910 : DMemory_769; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3935 = EXMEMop == 7'h23 ? _GEN_2911 : DMemory_770; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3936 = EXMEMop == 7'h23 ? _GEN_2912 : DMemory_771; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3937 = EXMEMop == 7'h23 ? _GEN_2913 : DMemory_772; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3938 = EXMEMop == 7'h23 ? _GEN_2914 : DMemory_773; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3939 = EXMEMop == 7'h23 ? _GEN_2915 : DMemory_774; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3940 = EXMEMop == 7'h23 ? _GEN_2916 : DMemory_775; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3941 = EXMEMop == 7'h23 ? _GEN_2917 : DMemory_776; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3942 = EXMEMop == 7'h23 ? _GEN_2918 : DMemory_777; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3943 = EXMEMop == 7'h23 ? _GEN_2919 : DMemory_778; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3944 = EXMEMop == 7'h23 ? _GEN_2920 : DMemory_779; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3945 = EXMEMop == 7'h23 ? _GEN_2921 : DMemory_780; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3946 = EXMEMop == 7'h23 ? _GEN_2922 : DMemory_781; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3947 = EXMEMop == 7'h23 ? _GEN_2923 : DMemory_782; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3948 = EXMEMop == 7'h23 ? _GEN_2924 : DMemory_783; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3949 = EXMEMop == 7'h23 ? _GEN_2925 : DMemory_784; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3950 = EXMEMop == 7'h23 ? _GEN_2926 : DMemory_785; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3951 = EXMEMop == 7'h23 ? _GEN_2927 : DMemory_786; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3952 = EXMEMop == 7'h23 ? _GEN_2928 : DMemory_787; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3953 = EXMEMop == 7'h23 ? _GEN_2929 : DMemory_788; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3954 = EXMEMop == 7'h23 ? _GEN_2930 : DMemory_789; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3955 = EXMEMop == 7'h23 ? _GEN_2931 : DMemory_790; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3956 = EXMEMop == 7'h23 ? _GEN_2932 : DMemory_791; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3957 = EXMEMop == 7'h23 ? _GEN_2933 : DMemory_792; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3958 = EXMEMop == 7'h23 ? _GEN_2934 : DMemory_793; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3959 = EXMEMop == 7'h23 ? _GEN_2935 : DMemory_794; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3960 = EXMEMop == 7'h23 ? _GEN_2936 : DMemory_795; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3961 = EXMEMop == 7'h23 ? _GEN_2937 : DMemory_796; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3962 = EXMEMop == 7'h23 ? _GEN_2938 : DMemory_797; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3963 = EXMEMop == 7'h23 ? _GEN_2939 : DMemory_798; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3964 = EXMEMop == 7'h23 ? _GEN_2940 : DMemory_799; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3965 = EXMEMop == 7'h23 ? _GEN_2941 : DMemory_800; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3966 = EXMEMop == 7'h23 ? _GEN_2942 : DMemory_801; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3967 = EXMEMop == 7'h23 ? _GEN_2943 : DMemory_802; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3968 = EXMEMop == 7'h23 ? _GEN_2944 : DMemory_803; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3969 = EXMEMop == 7'h23 ? _GEN_2945 : DMemory_804; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3970 = EXMEMop == 7'h23 ? _GEN_2946 : DMemory_805; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3971 = EXMEMop == 7'h23 ? _GEN_2947 : DMemory_806; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3972 = EXMEMop == 7'h23 ? _GEN_2948 : DMemory_807; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3973 = EXMEMop == 7'h23 ? _GEN_2949 : DMemory_808; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3974 = EXMEMop == 7'h23 ? _GEN_2950 : DMemory_809; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3975 = EXMEMop == 7'h23 ? _GEN_2951 : DMemory_810; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3976 = EXMEMop == 7'h23 ? _GEN_2952 : DMemory_811; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3977 = EXMEMop == 7'h23 ? _GEN_2953 : DMemory_812; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3978 = EXMEMop == 7'h23 ? _GEN_2954 : DMemory_813; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3979 = EXMEMop == 7'h23 ? _GEN_2955 : DMemory_814; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3980 = EXMEMop == 7'h23 ? _GEN_2956 : DMemory_815; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3981 = EXMEMop == 7'h23 ? _GEN_2957 : DMemory_816; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3982 = EXMEMop == 7'h23 ? _GEN_2958 : DMemory_817; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3983 = EXMEMop == 7'h23 ? _GEN_2959 : DMemory_818; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3984 = EXMEMop == 7'h23 ? _GEN_2960 : DMemory_819; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3985 = EXMEMop == 7'h23 ? _GEN_2961 : DMemory_820; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3986 = EXMEMop == 7'h23 ? _GEN_2962 : DMemory_821; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3987 = EXMEMop == 7'h23 ? _GEN_2963 : DMemory_822; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3988 = EXMEMop == 7'h23 ? _GEN_2964 : DMemory_823; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3989 = EXMEMop == 7'h23 ? _GEN_2965 : DMemory_824; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3990 = EXMEMop == 7'h23 ? _GEN_2966 : DMemory_825; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3991 = EXMEMop == 7'h23 ? _GEN_2967 : DMemory_826; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3992 = EXMEMop == 7'h23 ? _GEN_2968 : DMemory_827; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3993 = EXMEMop == 7'h23 ? _GEN_2969 : DMemory_828; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3994 = EXMEMop == 7'h23 ? _GEN_2970 : DMemory_829; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3995 = EXMEMop == 7'h23 ? _GEN_2971 : DMemory_830; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3996 = EXMEMop == 7'h23 ? _GEN_2972 : DMemory_831; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3997 = EXMEMop == 7'h23 ? _GEN_2973 : DMemory_832; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3998 = EXMEMop == 7'h23 ? _GEN_2974 : DMemory_833; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_3999 = EXMEMop == 7'h23 ? _GEN_2975 : DMemory_834; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4000 = EXMEMop == 7'h23 ? _GEN_2976 : DMemory_835; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4001 = EXMEMop == 7'h23 ? _GEN_2977 : DMemory_836; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4002 = EXMEMop == 7'h23 ? _GEN_2978 : DMemory_837; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4003 = EXMEMop == 7'h23 ? _GEN_2979 : DMemory_838; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4004 = EXMEMop == 7'h23 ? _GEN_2980 : DMemory_839; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4005 = EXMEMop == 7'h23 ? _GEN_2981 : DMemory_840; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4006 = EXMEMop == 7'h23 ? _GEN_2982 : DMemory_841; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4007 = EXMEMop == 7'h23 ? _GEN_2983 : DMemory_842; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4008 = EXMEMop == 7'h23 ? _GEN_2984 : DMemory_843; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4009 = EXMEMop == 7'h23 ? _GEN_2985 : DMemory_844; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4010 = EXMEMop == 7'h23 ? _GEN_2986 : DMemory_845; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4011 = EXMEMop == 7'h23 ? _GEN_2987 : DMemory_846; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4012 = EXMEMop == 7'h23 ? _GEN_2988 : DMemory_847; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4013 = EXMEMop == 7'h23 ? _GEN_2989 : DMemory_848; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4014 = EXMEMop == 7'h23 ? _GEN_2990 : DMemory_849; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4015 = EXMEMop == 7'h23 ? _GEN_2991 : DMemory_850; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4016 = EXMEMop == 7'h23 ? _GEN_2992 : DMemory_851; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4017 = EXMEMop == 7'h23 ? _GEN_2993 : DMemory_852; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4018 = EXMEMop == 7'h23 ? _GEN_2994 : DMemory_853; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4019 = EXMEMop == 7'h23 ? _GEN_2995 : DMemory_854; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4020 = EXMEMop == 7'h23 ? _GEN_2996 : DMemory_855; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4021 = EXMEMop == 7'h23 ? _GEN_2997 : DMemory_856; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4022 = EXMEMop == 7'h23 ? _GEN_2998 : DMemory_857; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4023 = EXMEMop == 7'h23 ? _GEN_2999 : DMemory_858; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4024 = EXMEMop == 7'h23 ? _GEN_3000 : DMemory_859; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4025 = EXMEMop == 7'h23 ? _GEN_3001 : DMemory_860; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4026 = EXMEMop == 7'h23 ? _GEN_3002 : DMemory_861; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4027 = EXMEMop == 7'h23 ? _GEN_3003 : DMemory_862; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4028 = EXMEMop == 7'h23 ? _GEN_3004 : DMemory_863; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4029 = EXMEMop == 7'h23 ? _GEN_3005 : DMemory_864; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4030 = EXMEMop == 7'h23 ? _GEN_3006 : DMemory_865; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4031 = EXMEMop == 7'h23 ? _GEN_3007 : DMemory_866; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4032 = EXMEMop == 7'h23 ? _GEN_3008 : DMemory_867; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4033 = EXMEMop == 7'h23 ? _GEN_3009 : DMemory_868; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4034 = EXMEMop == 7'h23 ? _GEN_3010 : DMemory_869; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4035 = EXMEMop == 7'h23 ? _GEN_3011 : DMemory_870; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4036 = EXMEMop == 7'h23 ? _GEN_3012 : DMemory_871; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4037 = EXMEMop == 7'h23 ? _GEN_3013 : DMemory_872; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4038 = EXMEMop == 7'h23 ? _GEN_3014 : DMemory_873; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4039 = EXMEMop == 7'h23 ? _GEN_3015 : DMemory_874; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4040 = EXMEMop == 7'h23 ? _GEN_3016 : DMemory_875; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4041 = EXMEMop == 7'h23 ? _GEN_3017 : DMemory_876; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4042 = EXMEMop == 7'h23 ? _GEN_3018 : DMemory_877; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4043 = EXMEMop == 7'h23 ? _GEN_3019 : DMemory_878; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4044 = EXMEMop == 7'h23 ? _GEN_3020 : DMemory_879; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4045 = EXMEMop == 7'h23 ? _GEN_3021 : DMemory_880; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4046 = EXMEMop == 7'h23 ? _GEN_3022 : DMemory_881; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4047 = EXMEMop == 7'h23 ? _GEN_3023 : DMemory_882; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4048 = EXMEMop == 7'h23 ? _GEN_3024 : DMemory_883; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4049 = EXMEMop == 7'h23 ? _GEN_3025 : DMemory_884; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4050 = EXMEMop == 7'h23 ? _GEN_3026 : DMemory_885; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4051 = EXMEMop == 7'h23 ? _GEN_3027 : DMemory_886; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4052 = EXMEMop == 7'h23 ? _GEN_3028 : DMemory_887; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4053 = EXMEMop == 7'h23 ? _GEN_3029 : DMemory_888; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4054 = EXMEMop == 7'h23 ? _GEN_3030 : DMemory_889; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4055 = EXMEMop == 7'h23 ? _GEN_3031 : DMemory_890; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4056 = EXMEMop == 7'h23 ? _GEN_3032 : DMemory_891; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4057 = EXMEMop == 7'h23 ? _GEN_3033 : DMemory_892; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4058 = EXMEMop == 7'h23 ? _GEN_3034 : DMemory_893; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4059 = EXMEMop == 7'h23 ? _GEN_3035 : DMemory_894; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4060 = EXMEMop == 7'h23 ? _GEN_3036 : DMemory_895; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4061 = EXMEMop == 7'h23 ? _GEN_3037 : DMemory_896; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4062 = EXMEMop == 7'h23 ? _GEN_3038 : DMemory_897; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4063 = EXMEMop == 7'h23 ? _GEN_3039 : DMemory_898; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4064 = EXMEMop == 7'h23 ? _GEN_3040 : DMemory_899; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4065 = EXMEMop == 7'h23 ? _GEN_3041 : DMemory_900; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4066 = EXMEMop == 7'h23 ? _GEN_3042 : DMemory_901; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4067 = EXMEMop == 7'h23 ? _GEN_3043 : DMemory_902; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4068 = EXMEMop == 7'h23 ? _GEN_3044 : DMemory_903; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4069 = EXMEMop == 7'h23 ? _GEN_3045 : DMemory_904; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4070 = EXMEMop == 7'h23 ? _GEN_3046 : DMemory_905; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4071 = EXMEMop == 7'h23 ? _GEN_3047 : DMemory_906; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4072 = EXMEMop == 7'h23 ? _GEN_3048 : DMemory_907; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4073 = EXMEMop == 7'h23 ? _GEN_3049 : DMemory_908; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4074 = EXMEMop == 7'h23 ? _GEN_3050 : DMemory_909; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4075 = EXMEMop == 7'h23 ? _GEN_3051 : DMemory_910; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4076 = EXMEMop == 7'h23 ? _GEN_3052 : DMemory_911; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4077 = EXMEMop == 7'h23 ? _GEN_3053 : DMemory_912; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4078 = EXMEMop == 7'h23 ? _GEN_3054 : DMemory_913; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4079 = EXMEMop == 7'h23 ? _GEN_3055 : DMemory_914; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4080 = EXMEMop == 7'h23 ? _GEN_3056 : DMemory_915; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4081 = EXMEMop == 7'h23 ? _GEN_3057 : DMemory_916; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4082 = EXMEMop == 7'h23 ? _GEN_3058 : DMemory_917; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4083 = EXMEMop == 7'h23 ? _GEN_3059 : DMemory_918; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4084 = EXMEMop == 7'h23 ? _GEN_3060 : DMemory_919; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4085 = EXMEMop == 7'h23 ? _GEN_3061 : DMemory_920; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4086 = EXMEMop == 7'h23 ? _GEN_3062 : DMemory_921; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4087 = EXMEMop == 7'h23 ? _GEN_3063 : DMemory_922; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4088 = EXMEMop == 7'h23 ? _GEN_3064 : DMemory_923; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4089 = EXMEMop == 7'h23 ? _GEN_3065 : DMemory_924; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4090 = EXMEMop == 7'h23 ? _GEN_3066 : DMemory_925; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4091 = EXMEMop == 7'h23 ? _GEN_3067 : DMemory_926; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4092 = EXMEMop == 7'h23 ? _GEN_3068 : DMemory_927; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4093 = EXMEMop == 7'h23 ? _GEN_3069 : DMemory_928; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4094 = EXMEMop == 7'h23 ? _GEN_3070 : DMemory_929; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4095 = EXMEMop == 7'h23 ? _GEN_3071 : DMemory_930; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4096 = EXMEMop == 7'h23 ? _GEN_3072 : DMemory_931; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4097 = EXMEMop == 7'h23 ? _GEN_3073 : DMemory_932; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4098 = EXMEMop == 7'h23 ? _GEN_3074 : DMemory_933; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4099 = EXMEMop == 7'h23 ? _GEN_3075 : DMemory_934; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4100 = EXMEMop == 7'h23 ? _GEN_3076 : DMemory_935; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4101 = EXMEMop == 7'h23 ? _GEN_3077 : DMemory_936; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4102 = EXMEMop == 7'h23 ? _GEN_3078 : DMemory_937; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4103 = EXMEMop == 7'h23 ? _GEN_3079 : DMemory_938; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4104 = EXMEMop == 7'h23 ? _GEN_3080 : DMemory_939; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4105 = EXMEMop == 7'h23 ? _GEN_3081 : DMemory_940; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4106 = EXMEMop == 7'h23 ? _GEN_3082 : DMemory_941; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4107 = EXMEMop == 7'h23 ? _GEN_3083 : DMemory_942; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4108 = EXMEMop == 7'h23 ? _GEN_3084 : DMemory_943; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4109 = EXMEMop == 7'h23 ? _GEN_3085 : DMemory_944; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4110 = EXMEMop == 7'h23 ? _GEN_3086 : DMemory_945; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4111 = EXMEMop == 7'h23 ? _GEN_3087 : DMemory_946; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4112 = EXMEMop == 7'h23 ? _GEN_3088 : DMemory_947; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4113 = EXMEMop == 7'h23 ? _GEN_3089 : DMemory_948; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4114 = EXMEMop == 7'h23 ? _GEN_3090 : DMemory_949; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4115 = EXMEMop == 7'h23 ? _GEN_3091 : DMemory_950; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4116 = EXMEMop == 7'h23 ? _GEN_3092 : DMemory_951; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4117 = EXMEMop == 7'h23 ? _GEN_3093 : DMemory_952; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4118 = EXMEMop == 7'h23 ? _GEN_3094 : DMemory_953; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4119 = EXMEMop == 7'h23 ? _GEN_3095 : DMemory_954; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4120 = EXMEMop == 7'h23 ? _GEN_3096 : DMemory_955; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4121 = EXMEMop == 7'h23 ? _GEN_3097 : DMemory_956; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4122 = EXMEMop == 7'h23 ? _GEN_3098 : DMemory_957; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4123 = EXMEMop == 7'h23 ? _GEN_3099 : DMemory_958; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4124 = EXMEMop == 7'h23 ? _GEN_3100 : DMemory_959; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4125 = EXMEMop == 7'h23 ? _GEN_3101 : DMemory_960; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4126 = EXMEMop == 7'h23 ? _GEN_3102 : DMemory_961; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4127 = EXMEMop == 7'h23 ? _GEN_3103 : DMemory_962; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4128 = EXMEMop == 7'h23 ? _GEN_3104 : DMemory_963; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4129 = EXMEMop == 7'h23 ? _GEN_3105 : DMemory_964; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4130 = EXMEMop == 7'h23 ? _GEN_3106 : DMemory_965; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4131 = EXMEMop == 7'h23 ? _GEN_3107 : DMemory_966; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4132 = EXMEMop == 7'h23 ? _GEN_3108 : DMemory_967; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4133 = EXMEMop == 7'h23 ? _GEN_3109 : DMemory_968; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4134 = EXMEMop == 7'h23 ? _GEN_3110 : DMemory_969; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4135 = EXMEMop == 7'h23 ? _GEN_3111 : DMemory_970; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4136 = EXMEMop == 7'h23 ? _GEN_3112 : DMemory_971; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4137 = EXMEMop == 7'h23 ? _GEN_3113 : DMemory_972; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4138 = EXMEMop == 7'h23 ? _GEN_3114 : DMemory_973; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4139 = EXMEMop == 7'h23 ? _GEN_3115 : DMemory_974; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4140 = EXMEMop == 7'h23 ? _GEN_3116 : DMemory_975; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4141 = EXMEMop == 7'h23 ? _GEN_3117 : DMemory_976; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4142 = EXMEMop == 7'h23 ? _GEN_3118 : DMemory_977; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4143 = EXMEMop == 7'h23 ? _GEN_3119 : DMemory_978; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4144 = EXMEMop == 7'h23 ? _GEN_3120 : DMemory_979; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4145 = EXMEMop == 7'h23 ? _GEN_3121 : DMemory_980; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4146 = EXMEMop == 7'h23 ? _GEN_3122 : DMemory_981; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4147 = EXMEMop == 7'h23 ? _GEN_3123 : DMemory_982; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4148 = EXMEMop == 7'h23 ? _GEN_3124 : DMemory_983; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4149 = EXMEMop == 7'h23 ? _GEN_3125 : DMemory_984; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4150 = EXMEMop == 7'h23 ? _GEN_3126 : DMemory_985; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4151 = EXMEMop == 7'h23 ? _GEN_3127 : DMemory_986; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4152 = EXMEMop == 7'h23 ? _GEN_3128 : DMemory_987; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4153 = EXMEMop == 7'h23 ? _GEN_3129 : DMemory_988; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4154 = EXMEMop == 7'h23 ? _GEN_3130 : DMemory_989; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4155 = EXMEMop == 7'h23 ? _GEN_3131 : DMemory_990; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4156 = EXMEMop == 7'h23 ? _GEN_3132 : DMemory_991; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4157 = EXMEMop == 7'h23 ? _GEN_3133 : DMemory_992; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4158 = EXMEMop == 7'h23 ? _GEN_3134 : DMemory_993; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4159 = EXMEMop == 7'h23 ? _GEN_3135 : DMemory_994; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4160 = EXMEMop == 7'h23 ? _GEN_3136 : DMemory_995; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4161 = EXMEMop == 7'h23 ? _GEN_3137 : DMemory_996; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4162 = EXMEMop == 7'h23 ? _GEN_3138 : DMemory_997; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4163 = EXMEMop == 7'h23 ? _GEN_3139 : DMemory_998; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4164 = EXMEMop == 7'h23 ? _GEN_3140 : DMemory_999; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4165 = EXMEMop == 7'h23 ? _GEN_3141 : DMemory_1000; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4166 = EXMEMop == 7'h23 ? _GEN_3142 : DMemory_1001; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4167 = EXMEMop == 7'h23 ? _GEN_3143 : DMemory_1002; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4168 = EXMEMop == 7'h23 ? _GEN_3144 : DMemory_1003; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4169 = EXMEMop == 7'h23 ? _GEN_3145 : DMemory_1004; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4170 = EXMEMop == 7'h23 ? _GEN_3146 : DMemory_1005; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4171 = EXMEMop == 7'h23 ? _GEN_3147 : DMemory_1006; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4172 = EXMEMop == 7'h23 ? _GEN_3148 : DMemory_1007; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4173 = EXMEMop == 7'h23 ? _GEN_3149 : DMemory_1008; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4174 = EXMEMop == 7'h23 ? _GEN_3150 : DMemory_1009; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4175 = EXMEMop == 7'h23 ? _GEN_3151 : DMemory_1010; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4176 = EXMEMop == 7'h23 ? _GEN_3152 : DMemory_1011; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4177 = EXMEMop == 7'h23 ? _GEN_3153 : DMemory_1012; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4178 = EXMEMop == 7'h23 ? _GEN_3154 : DMemory_1013; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4179 = EXMEMop == 7'h23 ? _GEN_3155 : DMemory_1014; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4180 = EXMEMop == 7'h23 ? _GEN_3156 : DMemory_1015; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4181 = EXMEMop == 7'h23 ? _GEN_3157 : DMemory_1016; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4182 = EXMEMop == 7'h23 ? _GEN_3158 : DMemory_1017; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4183 = EXMEMop == 7'h23 ? _GEN_3159 : DMemory_1018; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4184 = EXMEMop == 7'h23 ? _GEN_3160 : DMemory_1019; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4185 = EXMEMop == 7'h23 ? _GEN_3161 : DMemory_1020; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4186 = EXMEMop == 7'h23 ? _GEN_3162 : DMemory_1021; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4187 = EXMEMop == 7'h23 ? _GEN_3163 : DMemory_1022; // @[cpu.scala 220:32 69:24]
  wire [31:0] _GEN_4188 = EXMEMop == 7'h23 ? _GEN_3164 : DMemory_1023; // @[cpu.scala 220:32 69:24]
  assign io_rvfi_regs_0 = Regs_0; // @[cpu.scala 237:16]
  assign io_rvfi_regs_1 = Regs_1; // @[cpu.scala 237:16]
  assign io_rvfi_regs_2 = Regs_2; // @[cpu.scala 237:16]
  assign io_rvfi_regs_3 = Regs_3; // @[cpu.scala 237:16]
  assign io_rvfi_regs_4 = Regs_4; // @[cpu.scala 237:16]
  assign io_rvfi_regs_5 = Regs_5; // @[cpu.scala 237:16]
  assign io_rvfi_regs_6 = Regs_6; // @[cpu.scala 237:16]
  assign io_rvfi_regs_7 = Regs_7; // @[cpu.scala 237:16]
  assign io_rvfi_regs_8 = Regs_8; // @[cpu.scala 237:16]
  assign io_rvfi_regs_9 = Regs_9; // @[cpu.scala 237:16]
  assign io_rvfi_regs_10 = Regs_10; // @[cpu.scala 237:16]
  assign io_rvfi_regs_11 = Regs_11; // @[cpu.scala 237:16]
  assign io_rvfi_regs_12 = Regs_12; // @[cpu.scala 237:16]
  assign io_rvfi_regs_13 = Regs_13; // @[cpu.scala 237:16]
  assign io_rvfi_regs_14 = Regs_14; // @[cpu.scala 237:16]
  assign io_rvfi_regs_15 = Regs_15; // @[cpu.scala 237:16]
  assign io_rvfi_regs_16 = Regs_16; // @[cpu.scala 237:16]
  assign io_rvfi_regs_17 = Regs_17; // @[cpu.scala 237:16]
  assign io_rvfi_regs_18 = Regs_18; // @[cpu.scala 237:16]
  assign io_rvfi_regs_19 = Regs_19; // @[cpu.scala 237:16]
  assign io_rvfi_regs_20 = Regs_20; // @[cpu.scala 237:16]
  assign io_rvfi_regs_21 = Regs_21; // @[cpu.scala 237:16]
  assign io_rvfi_regs_22 = Regs_22; // @[cpu.scala 237:16]
  assign io_rvfi_regs_23 = Regs_23; // @[cpu.scala 237:16]
  assign io_rvfi_regs_24 = Regs_24; // @[cpu.scala 237:16]
  assign io_rvfi_regs_25 = Regs_25; // @[cpu.scala 237:16]
  assign io_rvfi_regs_26 = Regs_26; // @[cpu.scala 237:16]
  assign io_rvfi_regs_27 = Regs_27; // @[cpu.scala 237:16]
  assign io_rvfi_regs_28 = Regs_28; // @[cpu.scala 237:16]
  assign io_rvfi_regs_29 = Regs_29; // @[cpu.scala 237:16]
  assign io_rvfi_regs_30 = Regs_30; // @[cpu.scala 237:16]
  assign io_rvfi_regs_31 = Regs_31; // @[cpu.scala 237:16]
  always @(posedge clock) begin
    if (reset) begin // @[cpu.scala 64:19]
      PC <= 64'h0; // @[cpu.scala 64:19]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (~stall) begin // @[cpu.scala 137:27]
        if (~takeBranch) begin // @[cpu.scala 138:34]
          PC <= _PC_T_1; // @[cpu.scala 142:12]
        end else begin
          PC <= branchTarget; // @[cpu.scala 158:12]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_0 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h0 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_0 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_1 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h1 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_1 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_2 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h2 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_2 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_3 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h3 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_3 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_4 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h4 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_4 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_5 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h5 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_5 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_6 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h6 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_6 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_7 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h7 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_7 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_8 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h8 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_8 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_9 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h9 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_9 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_10 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'ha == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_10 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_11 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'hb == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_11 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_12 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'hc == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_12 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_13 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'hd == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_13 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_14 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'he == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_14 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_15 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'hf == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_15 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_16 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h10 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_16 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_17 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h11 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_17 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_18 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h12 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_18 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_19 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h13 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_19 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_20 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h14 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_20 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_21 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h15 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_21 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_22 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h16 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_22 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_23 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h17 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_23 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_24 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h18 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_24 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_25 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h19 == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_25 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_26 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h1a == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_26 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_27 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h1b == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_27 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_28 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h1c == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_28 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_29 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h1d == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_29 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_30 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h1e == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_30 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 65:21]
      Regs_31 <= 64'h0; // @[cpu.scala 65:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 230:74]
        if (5'h1f == MEMWBrd) begin // @[cpu.scala 231:21]
          Regs_31 <= MEMWBValue; // @[cpu.scala 231:21]
        end
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (~stall) begin // @[cpu.scala 137:27]
        if (bypassAFromEX) begin // @[cpu.scala 164:27]
          IDEXA <= _A_T_1; // @[cpu.scala 166:11]
        end else if (bypassAFromMEM) begin // @[cpu.scala 167:34]
          IDEXA <= EXMEMALUOut; // @[cpu.scala 169:11]
        end else begin
          IDEXA <= _GEN_1061;
        end
      end else begin
        IDEXA <= 64'h0;
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (~stall) begin // @[cpu.scala 137:27]
        if (bypassBFromEX) begin // @[cpu.scala 177:27]
          IDEXB <= _B_T_1; // @[cpu.scala 179:11]
        end else if (bypassBFromMEM) begin // @[cpu.scala 180:34]
          IDEXB <= EXMEMALUOut; // @[cpu.scala 182:11]
        end else begin
          IDEXB <= _GEN_1099;
        end
      end else begin
        IDEXB <= 64'h0;
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      EXMEMB <= IDEXB; // @[cpu.scala 213:12]
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (_stall_T_9) begin // @[cpu.scala 198:25]
        EXMEMALUOut <= _EXMEMALUOut_T_6; // @[cpu.scala 199:19]
      end else if (IDEXop == 7'h23) begin // @[cpu.scala 200:31]
        EXMEMALUOut <= _EXMEMALUOut_T_15; // @[cpu.scala 201:19]
      end else if (_bypassAFromEX_T_3) begin // @[cpu.scala 205:34]
        EXMEMALUOut <= _A_T_1; // @[cpu.scala 208:19]
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (_bypassAFromMEM_T_3) begin // @[cpu.scala 216:29]
        MEMWBValue <= EXMEMALUOut; // @[cpu.scala 217:18]
      end else if (_stall_T) begin // @[cpu.scala 218:32]
        MEMWBValue <= {{32'd0}, _GEN_2140}; // @[cpu.scala 219:18]
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_0 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_0 <= _GEN_3165;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1 <= _GEN_3166;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_2 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_2 <= _GEN_3167;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_3 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_3 <= _GEN_3168;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_4 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_4 <= _GEN_3169;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_5 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_5 <= _GEN_3170;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_6 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_6 <= _GEN_3171;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_7 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_7 <= _GEN_3172;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_8 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_8 <= _GEN_3173;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_9 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_9 <= _GEN_3174;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_10 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_10 <= _GEN_3175;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_11 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_11 <= _GEN_3176;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_12 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_12 <= _GEN_3177;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_13 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_13 <= _GEN_3178;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_14 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_14 <= _GEN_3179;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_15 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_15 <= _GEN_3180;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_16 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_16 <= _GEN_3181;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_17 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_17 <= _GEN_3182;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_18 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_18 <= _GEN_3183;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_19 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_19 <= _GEN_3184;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_20 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_20 <= _GEN_3185;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_21 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_21 <= _GEN_3186;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_22 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_22 <= _GEN_3187;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_23 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_23 <= _GEN_3188;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_24 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_24 <= _GEN_3189;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_25 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_25 <= _GEN_3190;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_26 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_26 <= _GEN_3191;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_27 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_27 <= _GEN_3192;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_28 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_28 <= _GEN_3193;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_29 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_29 <= _GEN_3194;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_30 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_30 <= _GEN_3195;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_31 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_31 <= _GEN_3196;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_32 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_32 <= _GEN_3197;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_33 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_33 <= _GEN_3198;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_34 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_34 <= _GEN_3199;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_35 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_35 <= _GEN_3200;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_36 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_36 <= _GEN_3201;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_37 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_37 <= _GEN_3202;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_38 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_38 <= _GEN_3203;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_39 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_39 <= _GEN_3204;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_40 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_40 <= _GEN_3205;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_41 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_41 <= _GEN_3206;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_42 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_42 <= _GEN_3207;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_43 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_43 <= _GEN_3208;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_44 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_44 <= _GEN_3209;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_45 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_45 <= _GEN_3210;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_46 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_46 <= _GEN_3211;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_47 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_47 <= _GEN_3212;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_48 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_48 <= _GEN_3213;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_49 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_49 <= _GEN_3214;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_50 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_50 <= _GEN_3215;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_51 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_51 <= _GEN_3216;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_52 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_52 <= _GEN_3217;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_53 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_53 <= _GEN_3218;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_54 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_54 <= _GEN_3219;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_55 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_55 <= _GEN_3220;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_56 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_56 <= _GEN_3221;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_57 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_57 <= _GEN_3222;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_58 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_58 <= _GEN_3223;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_59 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_59 <= _GEN_3224;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_60 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_60 <= _GEN_3225;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_61 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_61 <= _GEN_3226;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_62 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_62 <= _GEN_3227;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_63 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_63 <= _GEN_3228;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_64 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_64 <= _GEN_3229;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_65 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_65 <= _GEN_3230;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_66 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_66 <= _GEN_3231;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_67 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_67 <= _GEN_3232;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_68 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_68 <= _GEN_3233;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_69 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_69 <= _GEN_3234;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_70 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_70 <= _GEN_3235;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_71 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_71 <= _GEN_3236;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_72 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_72 <= _GEN_3237;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_73 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_73 <= _GEN_3238;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_74 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_74 <= _GEN_3239;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_75 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_75 <= _GEN_3240;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_76 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_76 <= _GEN_3241;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_77 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_77 <= _GEN_3242;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_78 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_78 <= _GEN_3243;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_79 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_79 <= _GEN_3244;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_80 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_80 <= _GEN_3245;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_81 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_81 <= _GEN_3246;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_82 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_82 <= _GEN_3247;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_83 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_83 <= _GEN_3248;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_84 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_84 <= _GEN_3249;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_85 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_85 <= _GEN_3250;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_86 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_86 <= _GEN_3251;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_87 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_87 <= _GEN_3252;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_88 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_88 <= _GEN_3253;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_89 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_89 <= _GEN_3254;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_90 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_90 <= _GEN_3255;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_91 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_91 <= _GEN_3256;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_92 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_92 <= _GEN_3257;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_93 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_93 <= _GEN_3258;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_94 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_94 <= _GEN_3259;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_95 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_95 <= _GEN_3260;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_96 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_96 <= _GEN_3261;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_97 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_97 <= _GEN_3262;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_98 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_98 <= _GEN_3263;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_99 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_99 <= _GEN_3264;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_100 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_100 <= _GEN_3265;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_101 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_101 <= _GEN_3266;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_102 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_102 <= _GEN_3267;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_103 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_103 <= _GEN_3268;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_104 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_104 <= _GEN_3269;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_105 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_105 <= _GEN_3270;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_106 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_106 <= _GEN_3271;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_107 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_107 <= _GEN_3272;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_108 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_108 <= _GEN_3273;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_109 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_109 <= _GEN_3274;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_110 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_110 <= _GEN_3275;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_111 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_111 <= _GEN_3276;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_112 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_112 <= _GEN_3277;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_113 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_113 <= _GEN_3278;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_114 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_114 <= _GEN_3279;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_115 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_115 <= _GEN_3280;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_116 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_116 <= _GEN_3281;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_117 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_117 <= _GEN_3282;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_118 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_118 <= _GEN_3283;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_119 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_119 <= _GEN_3284;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_120 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_120 <= _GEN_3285;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_121 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_121 <= _GEN_3286;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_122 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_122 <= _GEN_3287;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_123 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_123 <= _GEN_3288;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_124 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_124 <= _GEN_3289;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_125 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_125 <= _GEN_3290;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_126 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_126 <= _GEN_3291;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_127 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_127 <= _GEN_3292;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_128 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_128 <= _GEN_3293;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_129 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_129 <= _GEN_3294;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_130 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_130 <= _GEN_3295;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_131 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_131 <= _GEN_3296;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_132 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_132 <= _GEN_3297;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_133 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_133 <= _GEN_3298;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_134 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_134 <= _GEN_3299;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_135 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_135 <= _GEN_3300;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_136 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_136 <= _GEN_3301;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_137 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_137 <= _GEN_3302;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_138 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_138 <= _GEN_3303;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_139 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_139 <= _GEN_3304;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_140 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_140 <= _GEN_3305;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_141 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_141 <= _GEN_3306;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_142 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_142 <= _GEN_3307;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_143 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_143 <= _GEN_3308;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_144 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_144 <= _GEN_3309;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_145 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_145 <= _GEN_3310;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_146 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_146 <= _GEN_3311;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_147 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_147 <= _GEN_3312;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_148 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_148 <= _GEN_3313;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_149 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_149 <= _GEN_3314;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_150 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_150 <= _GEN_3315;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_151 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_151 <= _GEN_3316;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_152 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_152 <= _GEN_3317;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_153 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_153 <= _GEN_3318;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_154 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_154 <= _GEN_3319;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_155 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_155 <= _GEN_3320;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_156 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_156 <= _GEN_3321;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_157 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_157 <= _GEN_3322;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_158 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_158 <= _GEN_3323;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_159 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_159 <= _GEN_3324;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_160 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_160 <= _GEN_3325;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_161 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_161 <= _GEN_3326;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_162 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_162 <= _GEN_3327;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_163 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_163 <= _GEN_3328;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_164 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_164 <= _GEN_3329;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_165 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_165 <= _GEN_3330;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_166 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_166 <= _GEN_3331;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_167 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_167 <= _GEN_3332;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_168 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_168 <= _GEN_3333;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_169 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_169 <= _GEN_3334;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_170 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_170 <= _GEN_3335;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_171 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_171 <= _GEN_3336;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_172 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_172 <= _GEN_3337;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_173 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_173 <= _GEN_3338;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_174 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_174 <= _GEN_3339;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_175 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_175 <= _GEN_3340;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_176 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_176 <= _GEN_3341;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_177 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_177 <= _GEN_3342;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_178 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_178 <= _GEN_3343;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_179 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_179 <= _GEN_3344;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_180 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_180 <= _GEN_3345;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_181 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_181 <= _GEN_3346;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_182 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_182 <= _GEN_3347;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_183 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_183 <= _GEN_3348;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_184 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_184 <= _GEN_3349;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_185 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_185 <= _GEN_3350;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_186 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_186 <= _GEN_3351;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_187 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_187 <= _GEN_3352;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_188 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_188 <= _GEN_3353;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_189 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_189 <= _GEN_3354;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_190 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_190 <= _GEN_3355;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_191 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_191 <= _GEN_3356;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_192 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_192 <= _GEN_3357;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_193 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_193 <= _GEN_3358;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_194 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_194 <= _GEN_3359;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_195 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_195 <= _GEN_3360;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_196 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_196 <= _GEN_3361;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_197 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_197 <= _GEN_3362;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_198 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_198 <= _GEN_3363;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_199 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_199 <= _GEN_3364;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_200 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_200 <= _GEN_3365;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_201 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_201 <= _GEN_3366;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_202 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_202 <= _GEN_3367;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_203 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_203 <= _GEN_3368;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_204 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_204 <= _GEN_3369;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_205 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_205 <= _GEN_3370;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_206 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_206 <= _GEN_3371;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_207 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_207 <= _GEN_3372;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_208 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_208 <= _GEN_3373;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_209 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_209 <= _GEN_3374;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_210 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_210 <= _GEN_3375;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_211 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_211 <= _GEN_3376;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_212 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_212 <= _GEN_3377;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_213 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_213 <= _GEN_3378;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_214 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_214 <= _GEN_3379;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_215 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_215 <= _GEN_3380;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_216 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_216 <= _GEN_3381;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_217 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_217 <= _GEN_3382;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_218 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_218 <= _GEN_3383;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_219 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_219 <= _GEN_3384;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_220 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_220 <= _GEN_3385;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_221 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_221 <= _GEN_3386;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_222 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_222 <= _GEN_3387;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_223 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_223 <= _GEN_3388;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_224 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_224 <= _GEN_3389;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_225 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_225 <= _GEN_3390;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_226 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_226 <= _GEN_3391;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_227 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_227 <= _GEN_3392;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_228 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_228 <= _GEN_3393;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_229 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_229 <= _GEN_3394;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_230 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_230 <= _GEN_3395;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_231 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_231 <= _GEN_3396;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_232 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_232 <= _GEN_3397;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_233 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_233 <= _GEN_3398;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_234 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_234 <= _GEN_3399;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_235 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_235 <= _GEN_3400;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_236 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_236 <= _GEN_3401;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_237 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_237 <= _GEN_3402;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_238 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_238 <= _GEN_3403;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_239 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_239 <= _GEN_3404;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_240 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_240 <= _GEN_3405;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_241 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_241 <= _GEN_3406;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_242 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_242 <= _GEN_3407;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_243 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_243 <= _GEN_3408;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_244 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_244 <= _GEN_3409;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_245 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_245 <= _GEN_3410;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_246 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_246 <= _GEN_3411;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_247 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_247 <= _GEN_3412;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_248 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_248 <= _GEN_3413;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_249 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_249 <= _GEN_3414;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_250 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_250 <= _GEN_3415;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_251 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_251 <= _GEN_3416;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_252 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_252 <= _GEN_3417;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_253 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_253 <= _GEN_3418;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_254 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_254 <= _GEN_3419;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_255 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_255 <= _GEN_3420;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_256 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_256 <= _GEN_3421;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_257 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_257 <= _GEN_3422;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_258 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_258 <= _GEN_3423;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_259 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_259 <= _GEN_3424;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_260 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_260 <= _GEN_3425;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_261 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_261 <= _GEN_3426;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_262 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_262 <= _GEN_3427;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_263 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_263 <= _GEN_3428;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_264 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_264 <= _GEN_3429;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_265 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_265 <= _GEN_3430;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_266 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_266 <= _GEN_3431;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_267 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_267 <= _GEN_3432;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_268 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_268 <= _GEN_3433;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_269 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_269 <= _GEN_3434;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_270 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_270 <= _GEN_3435;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_271 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_271 <= _GEN_3436;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_272 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_272 <= _GEN_3437;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_273 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_273 <= _GEN_3438;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_274 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_274 <= _GEN_3439;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_275 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_275 <= _GEN_3440;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_276 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_276 <= _GEN_3441;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_277 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_277 <= _GEN_3442;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_278 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_278 <= _GEN_3443;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_279 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_279 <= _GEN_3444;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_280 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_280 <= _GEN_3445;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_281 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_281 <= _GEN_3446;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_282 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_282 <= _GEN_3447;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_283 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_283 <= _GEN_3448;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_284 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_284 <= _GEN_3449;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_285 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_285 <= _GEN_3450;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_286 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_286 <= _GEN_3451;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_287 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_287 <= _GEN_3452;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_288 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_288 <= _GEN_3453;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_289 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_289 <= _GEN_3454;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_290 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_290 <= _GEN_3455;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_291 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_291 <= _GEN_3456;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_292 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_292 <= _GEN_3457;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_293 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_293 <= _GEN_3458;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_294 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_294 <= _GEN_3459;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_295 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_295 <= _GEN_3460;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_296 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_296 <= _GEN_3461;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_297 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_297 <= _GEN_3462;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_298 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_298 <= _GEN_3463;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_299 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_299 <= _GEN_3464;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_300 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_300 <= _GEN_3465;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_301 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_301 <= _GEN_3466;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_302 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_302 <= _GEN_3467;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_303 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_303 <= _GEN_3468;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_304 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_304 <= _GEN_3469;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_305 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_305 <= _GEN_3470;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_306 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_306 <= _GEN_3471;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_307 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_307 <= _GEN_3472;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_308 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_308 <= _GEN_3473;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_309 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_309 <= _GEN_3474;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_310 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_310 <= _GEN_3475;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_311 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_311 <= _GEN_3476;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_312 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_312 <= _GEN_3477;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_313 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_313 <= _GEN_3478;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_314 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_314 <= _GEN_3479;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_315 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_315 <= _GEN_3480;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_316 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_316 <= _GEN_3481;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_317 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_317 <= _GEN_3482;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_318 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_318 <= _GEN_3483;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_319 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_319 <= _GEN_3484;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_320 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_320 <= _GEN_3485;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_321 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_321 <= _GEN_3486;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_322 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_322 <= _GEN_3487;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_323 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_323 <= _GEN_3488;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_324 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_324 <= _GEN_3489;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_325 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_325 <= _GEN_3490;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_326 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_326 <= _GEN_3491;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_327 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_327 <= _GEN_3492;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_328 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_328 <= _GEN_3493;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_329 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_329 <= _GEN_3494;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_330 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_330 <= _GEN_3495;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_331 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_331 <= _GEN_3496;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_332 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_332 <= _GEN_3497;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_333 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_333 <= _GEN_3498;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_334 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_334 <= _GEN_3499;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_335 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_335 <= _GEN_3500;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_336 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_336 <= _GEN_3501;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_337 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_337 <= _GEN_3502;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_338 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_338 <= _GEN_3503;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_339 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_339 <= _GEN_3504;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_340 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_340 <= _GEN_3505;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_341 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_341 <= _GEN_3506;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_342 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_342 <= _GEN_3507;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_343 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_343 <= _GEN_3508;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_344 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_344 <= _GEN_3509;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_345 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_345 <= _GEN_3510;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_346 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_346 <= _GEN_3511;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_347 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_347 <= _GEN_3512;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_348 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_348 <= _GEN_3513;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_349 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_349 <= _GEN_3514;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_350 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_350 <= _GEN_3515;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_351 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_351 <= _GEN_3516;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_352 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_352 <= _GEN_3517;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_353 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_353 <= _GEN_3518;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_354 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_354 <= _GEN_3519;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_355 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_355 <= _GEN_3520;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_356 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_356 <= _GEN_3521;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_357 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_357 <= _GEN_3522;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_358 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_358 <= _GEN_3523;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_359 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_359 <= _GEN_3524;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_360 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_360 <= _GEN_3525;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_361 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_361 <= _GEN_3526;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_362 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_362 <= _GEN_3527;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_363 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_363 <= _GEN_3528;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_364 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_364 <= _GEN_3529;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_365 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_365 <= _GEN_3530;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_366 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_366 <= _GEN_3531;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_367 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_367 <= _GEN_3532;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_368 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_368 <= _GEN_3533;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_369 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_369 <= _GEN_3534;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_370 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_370 <= _GEN_3535;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_371 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_371 <= _GEN_3536;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_372 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_372 <= _GEN_3537;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_373 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_373 <= _GEN_3538;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_374 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_374 <= _GEN_3539;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_375 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_375 <= _GEN_3540;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_376 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_376 <= _GEN_3541;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_377 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_377 <= _GEN_3542;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_378 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_378 <= _GEN_3543;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_379 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_379 <= _GEN_3544;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_380 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_380 <= _GEN_3545;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_381 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_381 <= _GEN_3546;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_382 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_382 <= _GEN_3547;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_383 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_383 <= _GEN_3548;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_384 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_384 <= _GEN_3549;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_385 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_385 <= _GEN_3550;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_386 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_386 <= _GEN_3551;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_387 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_387 <= _GEN_3552;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_388 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_388 <= _GEN_3553;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_389 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_389 <= _GEN_3554;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_390 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_390 <= _GEN_3555;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_391 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_391 <= _GEN_3556;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_392 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_392 <= _GEN_3557;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_393 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_393 <= _GEN_3558;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_394 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_394 <= _GEN_3559;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_395 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_395 <= _GEN_3560;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_396 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_396 <= _GEN_3561;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_397 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_397 <= _GEN_3562;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_398 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_398 <= _GEN_3563;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_399 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_399 <= _GEN_3564;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_400 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_400 <= _GEN_3565;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_401 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_401 <= _GEN_3566;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_402 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_402 <= _GEN_3567;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_403 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_403 <= _GEN_3568;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_404 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_404 <= _GEN_3569;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_405 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_405 <= _GEN_3570;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_406 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_406 <= _GEN_3571;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_407 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_407 <= _GEN_3572;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_408 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_408 <= _GEN_3573;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_409 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_409 <= _GEN_3574;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_410 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_410 <= _GEN_3575;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_411 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_411 <= _GEN_3576;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_412 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_412 <= _GEN_3577;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_413 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_413 <= _GEN_3578;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_414 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_414 <= _GEN_3579;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_415 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_415 <= _GEN_3580;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_416 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_416 <= _GEN_3581;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_417 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_417 <= _GEN_3582;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_418 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_418 <= _GEN_3583;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_419 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_419 <= _GEN_3584;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_420 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_420 <= _GEN_3585;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_421 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_421 <= _GEN_3586;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_422 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_422 <= _GEN_3587;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_423 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_423 <= _GEN_3588;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_424 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_424 <= _GEN_3589;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_425 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_425 <= _GEN_3590;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_426 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_426 <= _GEN_3591;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_427 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_427 <= _GEN_3592;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_428 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_428 <= _GEN_3593;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_429 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_429 <= _GEN_3594;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_430 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_430 <= _GEN_3595;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_431 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_431 <= _GEN_3596;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_432 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_432 <= _GEN_3597;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_433 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_433 <= _GEN_3598;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_434 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_434 <= _GEN_3599;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_435 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_435 <= _GEN_3600;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_436 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_436 <= _GEN_3601;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_437 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_437 <= _GEN_3602;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_438 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_438 <= _GEN_3603;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_439 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_439 <= _GEN_3604;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_440 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_440 <= _GEN_3605;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_441 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_441 <= _GEN_3606;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_442 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_442 <= _GEN_3607;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_443 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_443 <= _GEN_3608;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_444 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_444 <= _GEN_3609;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_445 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_445 <= _GEN_3610;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_446 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_446 <= _GEN_3611;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_447 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_447 <= _GEN_3612;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_448 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_448 <= _GEN_3613;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_449 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_449 <= _GEN_3614;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_450 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_450 <= _GEN_3615;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_451 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_451 <= _GEN_3616;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_452 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_452 <= _GEN_3617;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_453 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_453 <= _GEN_3618;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_454 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_454 <= _GEN_3619;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_455 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_455 <= _GEN_3620;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_456 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_456 <= _GEN_3621;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_457 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_457 <= _GEN_3622;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_458 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_458 <= _GEN_3623;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_459 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_459 <= _GEN_3624;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_460 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_460 <= _GEN_3625;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_461 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_461 <= _GEN_3626;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_462 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_462 <= _GEN_3627;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_463 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_463 <= _GEN_3628;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_464 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_464 <= _GEN_3629;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_465 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_465 <= _GEN_3630;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_466 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_466 <= _GEN_3631;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_467 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_467 <= _GEN_3632;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_468 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_468 <= _GEN_3633;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_469 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_469 <= _GEN_3634;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_470 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_470 <= _GEN_3635;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_471 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_471 <= _GEN_3636;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_472 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_472 <= _GEN_3637;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_473 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_473 <= _GEN_3638;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_474 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_474 <= _GEN_3639;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_475 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_475 <= _GEN_3640;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_476 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_476 <= _GEN_3641;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_477 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_477 <= _GEN_3642;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_478 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_478 <= _GEN_3643;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_479 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_479 <= _GEN_3644;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_480 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_480 <= _GEN_3645;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_481 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_481 <= _GEN_3646;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_482 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_482 <= _GEN_3647;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_483 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_483 <= _GEN_3648;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_484 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_484 <= _GEN_3649;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_485 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_485 <= _GEN_3650;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_486 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_486 <= _GEN_3651;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_487 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_487 <= _GEN_3652;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_488 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_488 <= _GEN_3653;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_489 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_489 <= _GEN_3654;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_490 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_490 <= _GEN_3655;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_491 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_491 <= _GEN_3656;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_492 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_492 <= _GEN_3657;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_493 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_493 <= _GEN_3658;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_494 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_494 <= _GEN_3659;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_495 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_495 <= _GEN_3660;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_496 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_496 <= _GEN_3661;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_497 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_497 <= _GEN_3662;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_498 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_498 <= _GEN_3663;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_499 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_499 <= _GEN_3664;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_500 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_500 <= _GEN_3665;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_501 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_501 <= _GEN_3666;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_502 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_502 <= _GEN_3667;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_503 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_503 <= _GEN_3668;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_504 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_504 <= _GEN_3669;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_505 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_505 <= _GEN_3670;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_506 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_506 <= _GEN_3671;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_507 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_507 <= _GEN_3672;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_508 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_508 <= _GEN_3673;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_509 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_509 <= _GEN_3674;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_510 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_510 <= _GEN_3675;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_511 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_511 <= _GEN_3676;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_512 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_512 <= _GEN_3677;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_513 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_513 <= _GEN_3678;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_514 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_514 <= _GEN_3679;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_515 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_515 <= _GEN_3680;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_516 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_516 <= _GEN_3681;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_517 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_517 <= _GEN_3682;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_518 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_518 <= _GEN_3683;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_519 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_519 <= _GEN_3684;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_520 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_520 <= _GEN_3685;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_521 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_521 <= _GEN_3686;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_522 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_522 <= _GEN_3687;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_523 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_523 <= _GEN_3688;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_524 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_524 <= _GEN_3689;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_525 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_525 <= _GEN_3690;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_526 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_526 <= _GEN_3691;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_527 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_527 <= _GEN_3692;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_528 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_528 <= _GEN_3693;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_529 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_529 <= _GEN_3694;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_530 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_530 <= _GEN_3695;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_531 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_531 <= _GEN_3696;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_532 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_532 <= _GEN_3697;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_533 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_533 <= _GEN_3698;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_534 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_534 <= _GEN_3699;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_535 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_535 <= _GEN_3700;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_536 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_536 <= _GEN_3701;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_537 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_537 <= _GEN_3702;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_538 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_538 <= _GEN_3703;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_539 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_539 <= _GEN_3704;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_540 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_540 <= _GEN_3705;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_541 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_541 <= _GEN_3706;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_542 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_542 <= _GEN_3707;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_543 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_543 <= _GEN_3708;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_544 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_544 <= _GEN_3709;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_545 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_545 <= _GEN_3710;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_546 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_546 <= _GEN_3711;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_547 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_547 <= _GEN_3712;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_548 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_548 <= _GEN_3713;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_549 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_549 <= _GEN_3714;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_550 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_550 <= _GEN_3715;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_551 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_551 <= _GEN_3716;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_552 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_552 <= _GEN_3717;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_553 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_553 <= _GEN_3718;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_554 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_554 <= _GEN_3719;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_555 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_555 <= _GEN_3720;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_556 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_556 <= _GEN_3721;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_557 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_557 <= _GEN_3722;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_558 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_558 <= _GEN_3723;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_559 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_559 <= _GEN_3724;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_560 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_560 <= _GEN_3725;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_561 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_561 <= _GEN_3726;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_562 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_562 <= _GEN_3727;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_563 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_563 <= _GEN_3728;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_564 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_564 <= _GEN_3729;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_565 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_565 <= _GEN_3730;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_566 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_566 <= _GEN_3731;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_567 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_567 <= _GEN_3732;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_568 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_568 <= _GEN_3733;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_569 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_569 <= _GEN_3734;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_570 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_570 <= _GEN_3735;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_571 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_571 <= _GEN_3736;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_572 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_572 <= _GEN_3737;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_573 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_573 <= _GEN_3738;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_574 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_574 <= _GEN_3739;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_575 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_575 <= _GEN_3740;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_576 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_576 <= _GEN_3741;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_577 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_577 <= _GEN_3742;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_578 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_578 <= _GEN_3743;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_579 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_579 <= _GEN_3744;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_580 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_580 <= _GEN_3745;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_581 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_581 <= _GEN_3746;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_582 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_582 <= _GEN_3747;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_583 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_583 <= _GEN_3748;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_584 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_584 <= _GEN_3749;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_585 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_585 <= _GEN_3750;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_586 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_586 <= _GEN_3751;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_587 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_587 <= _GEN_3752;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_588 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_588 <= _GEN_3753;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_589 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_589 <= _GEN_3754;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_590 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_590 <= _GEN_3755;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_591 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_591 <= _GEN_3756;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_592 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_592 <= _GEN_3757;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_593 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_593 <= _GEN_3758;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_594 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_594 <= _GEN_3759;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_595 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_595 <= _GEN_3760;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_596 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_596 <= _GEN_3761;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_597 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_597 <= _GEN_3762;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_598 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_598 <= _GEN_3763;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_599 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_599 <= _GEN_3764;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_600 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_600 <= _GEN_3765;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_601 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_601 <= _GEN_3766;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_602 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_602 <= _GEN_3767;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_603 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_603 <= _GEN_3768;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_604 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_604 <= _GEN_3769;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_605 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_605 <= _GEN_3770;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_606 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_606 <= _GEN_3771;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_607 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_607 <= _GEN_3772;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_608 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_608 <= _GEN_3773;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_609 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_609 <= _GEN_3774;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_610 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_610 <= _GEN_3775;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_611 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_611 <= _GEN_3776;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_612 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_612 <= _GEN_3777;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_613 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_613 <= _GEN_3778;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_614 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_614 <= _GEN_3779;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_615 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_615 <= _GEN_3780;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_616 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_616 <= _GEN_3781;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_617 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_617 <= _GEN_3782;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_618 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_618 <= _GEN_3783;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_619 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_619 <= _GEN_3784;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_620 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_620 <= _GEN_3785;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_621 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_621 <= _GEN_3786;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_622 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_622 <= _GEN_3787;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_623 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_623 <= _GEN_3788;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_624 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_624 <= _GEN_3789;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_625 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_625 <= _GEN_3790;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_626 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_626 <= _GEN_3791;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_627 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_627 <= _GEN_3792;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_628 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_628 <= _GEN_3793;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_629 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_629 <= _GEN_3794;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_630 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_630 <= _GEN_3795;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_631 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_631 <= _GEN_3796;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_632 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_632 <= _GEN_3797;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_633 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_633 <= _GEN_3798;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_634 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_634 <= _GEN_3799;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_635 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_635 <= _GEN_3800;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_636 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_636 <= _GEN_3801;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_637 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_637 <= _GEN_3802;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_638 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_638 <= _GEN_3803;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_639 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_639 <= _GEN_3804;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_640 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_640 <= _GEN_3805;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_641 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_641 <= _GEN_3806;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_642 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_642 <= _GEN_3807;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_643 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_643 <= _GEN_3808;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_644 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_644 <= _GEN_3809;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_645 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_645 <= _GEN_3810;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_646 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_646 <= _GEN_3811;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_647 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_647 <= _GEN_3812;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_648 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_648 <= _GEN_3813;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_649 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_649 <= _GEN_3814;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_650 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_650 <= _GEN_3815;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_651 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_651 <= _GEN_3816;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_652 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_652 <= _GEN_3817;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_653 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_653 <= _GEN_3818;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_654 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_654 <= _GEN_3819;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_655 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_655 <= _GEN_3820;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_656 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_656 <= _GEN_3821;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_657 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_657 <= _GEN_3822;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_658 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_658 <= _GEN_3823;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_659 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_659 <= _GEN_3824;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_660 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_660 <= _GEN_3825;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_661 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_661 <= _GEN_3826;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_662 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_662 <= _GEN_3827;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_663 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_663 <= _GEN_3828;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_664 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_664 <= _GEN_3829;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_665 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_665 <= _GEN_3830;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_666 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_666 <= _GEN_3831;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_667 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_667 <= _GEN_3832;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_668 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_668 <= _GEN_3833;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_669 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_669 <= _GEN_3834;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_670 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_670 <= _GEN_3835;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_671 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_671 <= _GEN_3836;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_672 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_672 <= _GEN_3837;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_673 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_673 <= _GEN_3838;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_674 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_674 <= _GEN_3839;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_675 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_675 <= _GEN_3840;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_676 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_676 <= _GEN_3841;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_677 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_677 <= _GEN_3842;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_678 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_678 <= _GEN_3843;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_679 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_679 <= _GEN_3844;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_680 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_680 <= _GEN_3845;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_681 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_681 <= _GEN_3846;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_682 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_682 <= _GEN_3847;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_683 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_683 <= _GEN_3848;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_684 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_684 <= _GEN_3849;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_685 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_685 <= _GEN_3850;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_686 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_686 <= _GEN_3851;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_687 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_687 <= _GEN_3852;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_688 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_688 <= _GEN_3853;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_689 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_689 <= _GEN_3854;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_690 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_690 <= _GEN_3855;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_691 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_691 <= _GEN_3856;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_692 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_692 <= _GEN_3857;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_693 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_693 <= _GEN_3858;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_694 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_694 <= _GEN_3859;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_695 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_695 <= _GEN_3860;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_696 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_696 <= _GEN_3861;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_697 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_697 <= _GEN_3862;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_698 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_698 <= _GEN_3863;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_699 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_699 <= _GEN_3864;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_700 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_700 <= _GEN_3865;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_701 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_701 <= _GEN_3866;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_702 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_702 <= _GEN_3867;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_703 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_703 <= _GEN_3868;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_704 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_704 <= _GEN_3869;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_705 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_705 <= _GEN_3870;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_706 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_706 <= _GEN_3871;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_707 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_707 <= _GEN_3872;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_708 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_708 <= _GEN_3873;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_709 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_709 <= _GEN_3874;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_710 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_710 <= _GEN_3875;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_711 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_711 <= _GEN_3876;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_712 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_712 <= _GEN_3877;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_713 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_713 <= _GEN_3878;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_714 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_714 <= _GEN_3879;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_715 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_715 <= _GEN_3880;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_716 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_716 <= _GEN_3881;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_717 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_717 <= _GEN_3882;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_718 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_718 <= _GEN_3883;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_719 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_719 <= _GEN_3884;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_720 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_720 <= _GEN_3885;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_721 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_721 <= _GEN_3886;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_722 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_722 <= _GEN_3887;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_723 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_723 <= _GEN_3888;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_724 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_724 <= _GEN_3889;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_725 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_725 <= _GEN_3890;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_726 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_726 <= _GEN_3891;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_727 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_727 <= _GEN_3892;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_728 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_728 <= _GEN_3893;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_729 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_729 <= _GEN_3894;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_730 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_730 <= _GEN_3895;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_731 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_731 <= _GEN_3896;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_732 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_732 <= _GEN_3897;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_733 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_733 <= _GEN_3898;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_734 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_734 <= _GEN_3899;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_735 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_735 <= _GEN_3900;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_736 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_736 <= _GEN_3901;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_737 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_737 <= _GEN_3902;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_738 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_738 <= _GEN_3903;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_739 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_739 <= _GEN_3904;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_740 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_740 <= _GEN_3905;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_741 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_741 <= _GEN_3906;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_742 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_742 <= _GEN_3907;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_743 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_743 <= _GEN_3908;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_744 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_744 <= _GEN_3909;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_745 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_745 <= _GEN_3910;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_746 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_746 <= _GEN_3911;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_747 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_747 <= _GEN_3912;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_748 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_748 <= _GEN_3913;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_749 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_749 <= _GEN_3914;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_750 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_750 <= _GEN_3915;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_751 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_751 <= _GEN_3916;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_752 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_752 <= _GEN_3917;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_753 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_753 <= _GEN_3918;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_754 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_754 <= _GEN_3919;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_755 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_755 <= _GEN_3920;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_756 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_756 <= _GEN_3921;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_757 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_757 <= _GEN_3922;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_758 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_758 <= _GEN_3923;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_759 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_759 <= _GEN_3924;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_760 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_760 <= _GEN_3925;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_761 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_761 <= _GEN_3926;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_762 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_762 <= _GEN_3927;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_763 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_763 <= _GEN_3928;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_764 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_764 <= _GEN_3929;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_765 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_765 <= _GEN_3930;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_766 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_766 <= _GEN_3931;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_767 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_767 <= _GEN_3932;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_768 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_768 <= _GEN_3933;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_769 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_769 <= _GEN_3934;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_770 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_770 <= _GEN_3935;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_771 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_771 <= _GEN_3936;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_772 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_772 <= _GEN_3937;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_773 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_773 <= _GEN_3938;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_774 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_774 <= _GEN_3939;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_775 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_775 <= _GEN_3940;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_776 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_776 <= _GEN_3941;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_777 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_777 <= _GEN_3942;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_778 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_778 <= _GEN_3943;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_779 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_779 <= _GEN_3944;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_780 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_780 <= _GEN_3945;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_781 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_781 <= _GEN_3946;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_782 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_782 <= _GEN_3947;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_783 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_783 <= _GEN_3948;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_784 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_784 <= _GEN_3949;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_785 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_785 <= _GEN_3950;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_786 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_786 <= _GEN_3951;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_787 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_787 <= _GEN_3952;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_788 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_788 <= _GEN_3953;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_789 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_789 <= _GEN_3954;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_790 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_790 <= _GEN_3955;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_791 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_791 <= _GEN_3956;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_792 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_792 <= _GEN_3957;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_793 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_793 <= _GEN_3958;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_794 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_794 <= _GEN_3959;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_795 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_795 <= _GEN_3960;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_796 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_796 <= _GEN_3961;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_797 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_797 <= _GEN_3962;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_798 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_798 <= _GEN_3963;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_799 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_799 <= _GEN_3964;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_800 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_800 <= _GEN_3965;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_801 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_801 <= _GEN_3966;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_802 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_802 <= _GEN_3967;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_803 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_803 <= _GEN_3968;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_804 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_804 <= _GEN_3969;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_805 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_805 <= _GEN_3970;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_806 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_806 <= _GEN_3971;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_807 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_807 <= _GEN_3972;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_808 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_808 <= _GEN_3973;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_809 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_809 <= _GEN_3974;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_810 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_810 <= _GEN_3975;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_811 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_811 <= _GEN_3976;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_812 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_812 <= _GEN_3977;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_813 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_813 <= _GEN_3978;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_814 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_814 <= _GEN_3979;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_815 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_815 <= _GEN_3980;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_816 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_816 <= _GEN_3981;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_817 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_817 <= _GEN_3982;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_818 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_818 <= _GEN_3983;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_819 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_819 <= _GEN_3984;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_820 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_820 <= _GEN_3985;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_821 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_821 <= _GEN_3986;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_822 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_822 <= _GEN_3987;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_823 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_823 <= _GEN_3988;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_824 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_824 <= _GEN_3989;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_825 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_825 <= _GEN_3990;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_826 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_826 <= _GEN_3991;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_827 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_827 <= _GEN_3992;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_828 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_828 <= _GEN_3993;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_829 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_829 <= _GEN_3994;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_830 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_830 <= _GEN_3995;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_831 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_831 <= _GEN_3996;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_832 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_832 <= _GEN_3997;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_833 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_833 <= _GEN_3998;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_834 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_834 <= _GEN_3999;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_835 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_835 <= _GEN_4000;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_836 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_836 <= _GEN_4001;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_837 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_837 <= _GEN_4002;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_838 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_838 <= _GEN_4003;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_839 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_839 <= _GEN_4004;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_840 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_840 <= _GEN_4005;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_841 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_841 <= _GEN_4006;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_842 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_842 <= _GEN_4007;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_843 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_843 <= _GEN_4008;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_844 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_844 <= _GEN_4009;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_845 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_845 <= _GEN_4010;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_846 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_846 <= _GEN_4011;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_847 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_847 <= _GEN_4012;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_848 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_848 <= _GEN_4013;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_849 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_849 <= _GEN_4014;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_850 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_850 <= _GEN_4015;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_851 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_851 <= _GEN_4016;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_852 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_852 <= _GEN_4017;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_853 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_853 <= _GEN_4018;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_854 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_854 <= _GEN_4019;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_855 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_855 <= _GEN_4020;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_856 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_856 <= _GEN_4021;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_857 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_857 <= _GEN_4022;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_858 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_858 <= _GEN_4023;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_859 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_859 <= _GEN_4024;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_860 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_860 <= _GEN_4025;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_861 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_861 <= _GEN_4026;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_862 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_862 <= _GEN_4027;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_863 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_863 <= _GEN_4028;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_864 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_864 <= _GEN_4029;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_865 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_865 <= _GEN_4030;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_866 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_866 <= _GEN_4031;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_867 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_867 <= _GEN_4032;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_868 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_868 <= _GEN_4033;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_869 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_869 <= _GEN_4034;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_870 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_870 <= _GEN_4035;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_871 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_871 <= _GEN_4036;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_872 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_872 <= _GEN_4037;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_873 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_873 <= _GEN_4038;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_874 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_874 <= _GEN_4039;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_875 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_875 <= _GEN_4040;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_876 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_876 <= _GEN_4041;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_877 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_877 <= _GEN_4042;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_878 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_878 <= _GEN_4043;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_879 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_879 <= _GEN_4044;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_880 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_880 <= _GEN_4045;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_881 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_881 <= _GEN_4046;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_882 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_882 <= _GEN_4047;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_883 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_883 <= _GEN_4048;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_884 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_884 <= _GEN_4049;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_885 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_885 <= _GEN_4050;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_886 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_886 <= _GEN_4051;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_887 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_887 <= _GEN_4052;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_888 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_888 <= _GEN_4053;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_889 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_889 <= _GEN_4054;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_890 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_890 <= _GEN_4055;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_891 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_891 <= _GEN_4056;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_892 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_892 <= _GEN_4057;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_893 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_893 <= _GEN_4058;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_894 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_894 <= _GEN_4059;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_895 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_895 <= _GEN_4060;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_896 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_896 <= _GEN_4061;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_897 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_897 <= _GEN_4062;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_898 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_898 <= _GEN_4063;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_899 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_899 <= _GEN_4064;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_900 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_900 <= _GEN_4065;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_901 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_901 <= _GEN_4066;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_902 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_902 <= _GEN_4067;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_903 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_903 <= _GEN_4068;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_904 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_904 <= _GEN_4069;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_905 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_905 <= _GEN_4070;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_906 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_906 <= _GEN_4071;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_907 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_907 <= _GEN_4072;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_908 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_908 <= _GEN_4073;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_909 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_909 <= _GEN_4074;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_910 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_910 <= _GEN_4075;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_911 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_911 <= _GEN_4076;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_912 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_912 <= _GEN_4077;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_913 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_913 <= _GEN_4078;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_914 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_914 <= _GEN_4079;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_915 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_915 <= _GEN_4080;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_916 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_916 <= _GEN_4081;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_917 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_917 <= _GEN_4082;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_918 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_918 <= _GEN_4083;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_919 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_919 <= _GEN_4084;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_920 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_920 <= _GEN_4085;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_921 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_921 <= _GEN_4086;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_922 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_922 <= _GEN_4087;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_923 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_923 <= _GEN_4088;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_924 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_924 <= _GEN_4089;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_925 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_925 <= _GEN_4090;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_926 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_926 <= _GEN_4091;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_927 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_927 <= _GEN_4092;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_928 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_928 <= _GEN_4093;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_929 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_929 <= _GEN_4094;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_930 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_930 <= _GEN_4095;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_931 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_931 <= _GEN_4096;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_932 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_932 <= _GEN_4097;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_933 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_933 <= _GEN_4098;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_934 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_934 <= _GEN_4099;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_935 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_935 <= _GEN_4100;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_936 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_936 <= _GEN_4101;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_937 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_937 <= _GEN_4102;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_938 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_938 <= _GEN_4103;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_939 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_939 <= _GEN_4104;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_940 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_940 <= _GEN_4105;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_941 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_941 <= _GEN_4106;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_942 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_942 <= _GEN_4107;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_943 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_943 <= _GEN_4108;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_944 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_944 <= _GEN_4109;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_945 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_945 <= _GEN_4110;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_946 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_946 <= _GEN_4111;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_947 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_947 <= _GEN_4112;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_948 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_948 <= _GEN_4113;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_949 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_949 <= _GEN_4114;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_950 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_950 <= _GEN_4115;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_951 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_951 <= _GEN_4116;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_952 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_952 <= _GEN_4117;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_953 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_953 <= _GEN_4118;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_954 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_954 <= _GEN_4119;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_955 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_955 <= _GEN_4120;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_956 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_956 <= _GEN_4121;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_957 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_957 <= _GEN_4122;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_958 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_958 <= _GEN_4123;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_959 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_959 <= _GEN_4124;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_960 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_960 <= _GEN_4125;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_961 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_961 <= _GEN_4126;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_962 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_962 <= _GEN_4127;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_963 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_963 <= _GEN_4128;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_964 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_964 <= _GEN_4129;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_965 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_965 <= _GEN_4130;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_966 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_966 <= _GEN_4131;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_967 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_967 <= _GEN_4132;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_968 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_968 <= _GEN_4133;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_969 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_969 <= _GEN_4134;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_970 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_970 <= _GEN_4135;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_971 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_971 <= _GEN_4136;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_972 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_972 <= _GEN_4137;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_973 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_973 <= _GEN_4138;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_974 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_974 <= _GEN_4139;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_975 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_975 <= _GEN_4140;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_976 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_976 <= _GEN_4141;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_977 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_977 <= _GEN_4142;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_978 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_978 <= _GEN_4143;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_979 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_979 <= _GEN_4144;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_980 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_980 <= _GEN_4145;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_981 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_981 <= _GEN_4146;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_982 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_982 <= _GEN_4147;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_983 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_983 <= _GEN_4148;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_984 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_984 <= _GEN_4149;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_985 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_985 <= _GEN_4150;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_986 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_986 <= _GEN_4151;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_987 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_987 <= _GEN_4152;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_988 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_988 <= _GEN_4153;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_989 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_989 <= _GEN_4154;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_990 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_990 <= _GEN_4155;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_991 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_991 <= _GEN_4156;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_992 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_992 <= _GEN_4157;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_993 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_993 <= _GEN_4158;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_994 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_994 <= _GEN_4159;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_995 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_995 <= _GEN_4160;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_996 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_996 <= _GEN_4161;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_997 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_997 <= _GEN_4162;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_998 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_998 <= _GEN_4163;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_999 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_999 <= _GEN_4164;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1000 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1000 <= _GEN_4165;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1001 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1001 <= _GEN_4166;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1002 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1002 <= _GEN_4167;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1003 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1003 <= _GEN_4168;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1004 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1004 <= _GEN_4169;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1005 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1005 <= _GEN_4170;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1006 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1006 <= _GEN_4171;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1007 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1007 <= _GEN_4172;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1008 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1008 <= _GEN_4173;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1009 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1009 <= _GEN_4174;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1010 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1010 <= _GEN_4175;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1011 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1011 <= _GEN_4176;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1012 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1012 <= _GEN_4177;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1013 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1013 <= _GEN_4178;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1014 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1014 <= _GEN_4179;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1015 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1015 <= _GEN_4180;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1016 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1016 <= _GEN_4181;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1017 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1017 <= _GEN_4182;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1018 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1018 <= _GEN_4183;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1019 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1019 <= _GEN_4184;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1020 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1020 <= _GEN_4185;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1021 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1021 <= _GEN_4186;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1022 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1022 <= _GEN_4187;
        end
      end
    end
    if (reset) begin // @[cpu.scala 69:24]
      DMemory_1023 <= 32'h0; // @[cpu.scala 69:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 216:29]
        if (!(_stall_T)) begin // @[cpu.scala 218:32]
          DMemory_1023 <= _GEN_4188;
        end
      end
    end
    if (reset) begin // @[cpu.scala 70:24]
      IMemory_0 <= 32'h13; // @[cpu.scala 70:24]
    end else if (io_rvfi_rst) begin // @[cpu.scala 80:21]
      IMemory_0 <= io_rvfi_insn_in_0; // @[cpu.scala 90:18]
    end
    if (reset) begin // @[cpu.scala 70:24]
      IMemory_1 <= 32'h13; // @[cpu.scala 70:24]
    end else if (io_rvfi_rst) begin // @[cpu.scala 80:21]
      IMemory_1 <= io_rvfi_insn_in_1; // @[cpu.scala 90:18]
    end
    if (reset) begin // @[cpu.scala 73:49]
      IFIDIR <= 32'h13; // @[cpu.scala 73:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (~stall) begin // @[cpu.scala 137:27]
        if (~takeBranch) begin // @[cpu.scala 138:34]
          IFIDIR <= _GEN_1023; // @[cpu.scala 141:16]
        end else begin
          IFIDIR <= 32'h13; // @[cpu.scala 145:16]
        end
      end
    end
    if (reset) begin // @[cpu.scala 73:49]
      IDEXIR <= 32'h13; // @[cpu.scala 73:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (~stall) begin // @[cpu.scala 137:27]
        IDEXIR <= IFIDIR; // @[cpu.scala 190:14]
      end else begin
        IDEXIR <= 32'h13; // @[cpu.scala 192:14]
      end
    end
    if (reset) begin // @[cpu.scala 73:49]
      EXMEMIR <= 32'h13; // @[cpu.scala 73:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      EXMEMIR <= IDEXIR; // @[cpu.scala 212:13]
    end
    if (reset) begin // @[cpu.scala 73:49]
      MEMWBIR <= 32'h13; // @[cpu.scala 73:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      MEMWBIR <= EXMEMIR; // @[cpu.scala 224:13]
    end
    if (reset) begin // @[cpu.scala 76:22]
      CurPC <= 64'h0; // @[cpu.scala 76:22]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 80:21]
      if (~stall) begin // @[cpu.scala 137:27]
        CurPC <= PC; // @[cpu.scala 161:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  PC = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  Regs_0 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  Regs_1 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  Regs_2 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  Regs_3 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  Regs_4 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  Regs_5 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  Regs_6 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  Regs_7 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  Regs_8 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  Regs_9 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  Regs_10 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  Regs_11 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  Regs_12 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  Regs_13 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  Regs_14 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  Regs_15 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  Regs_16 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  Regs_17 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  Regs_18 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  Regs_19 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  Regs_20 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  Regs_21 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  Regs_22 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  Regs_23 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  Regs_24 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  Regs_25 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  Regs_26 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  Regs_27 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  Regs_28 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  Regs_29 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  Regs_30 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  Regs_31 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  IDEXA = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  IDEXB = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  EXMEMB = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  EXMEMALUOut = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  MEMWBValue = _RAND_37[63:0];
  _RAND_38 = {1{`RANDOM}};
  DMemory_0 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  DMemory_1 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  DMemory_2 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  DMemory_3 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  DMemory_4 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  DMemory_5 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  DMemory_6 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  DMemory_7 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  DMemory_8 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  DMemory_9 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  DMemory_10 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  DMemory_11 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  DMemory_12 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  DMemory_13 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  DMemory_14 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  DMemory_15 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  DMemory_16 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  DMemory_17 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  DMemory_18 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  DMemory_19 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  DMemory_20 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  DMemory_21 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  DMemory_22 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  DMemory_23 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  DMemory_24 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  DMemory_25 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  DMemory_26 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  DMemory_27 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  DMemory_28 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  DMemory_29 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  DMemory_30 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  DMemory_31 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  DMemory_32 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  DMemory_33 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  DMemory_34 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  DMemory_35 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  DMemory_36 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  DMemory_37 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  DMemory_38 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  DMemory_39 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  DMemory_40 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  DMemory_41 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  DMemory_42 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  DMemory_43 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  DMemory_44 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  DMemory_45 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  DMemory_46 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  DMemory_47 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  DMemory_48 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  DMemory_49 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  DMemory_50 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  DMemory_51 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  DMemory_52 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  DMemory_53 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  DMemory_54 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  DMemory_55 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  DMemory_56 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  DMemory_57 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  DMemory_58 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  DMemory_59 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  DMemory_60 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  DMemory_61 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  DMemory_62 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  DMemory_63 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  DMemory_64 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  DMemory_65 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  DMemory_66 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  DMemory_67 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  DMemory_68 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  DMemory_69 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  DMemory_70 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  DMemory_71 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  DMemory_72 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  DMemory_73 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  DMemory_74 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  DMemory_75 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  DMemory_76 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  DMemory_77 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  DMemory_78 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  DMemory_79 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  DMemory_80 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  DMemory_81 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  DMemory_82 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  DMemory_83 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  DMemory_84 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  DMemory_85 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  DMemory_86 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  DMemory_87 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  DMemory_88 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  DMemory_89 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  DMemory_90 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  DMemory_91 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  DMemory_92 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  DMemory_93 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  DMemory_94 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  DMemory_95 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  DMemory_96 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  DMemory_97 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  DMemory_98 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  DMemory_99 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  DMemory_100 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  DMemory_101 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  DMemory_102 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  DMemory_103 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  DMemory_104 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  DMemory_105 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  DMemory_106 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  DMemory_107 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  DMemory_108 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  DMemory_109 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  DMemory_110 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  DMemory_111 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  DMemory_112 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  DMemory_113 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  DMemory_114 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  DMemory_115 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  DMemory_116 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  DMemory_117 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  DMemory_118 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  DMemory_119 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  DMemory_120 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  DMemory_121 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  DMemory_122 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  DMemory_123 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  DMemory_124 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  DMemory_125 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  DMemory_126 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  DMemory_127 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  DMemory_128 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  DMemory_129 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  DMemory_130 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  DMemory_131 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  DMemory_132 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  DMemory_133 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  DMemory_134 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  DMemory_135 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  DMemory_136 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  DMemory_137 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  DMemory_138 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  DMemory_139 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  DMemory_140 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  DMemory_141 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  DMemory_142 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  DMemory_143 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  DMemory_144 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  DMemory_145 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  DMemory_146 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  DMemory_147 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  DMemory_148 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  DMemory_149 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  DMemory_150 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  DMemory_151 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  DMemory_152 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  DMemory_153 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  DMemory_154 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  DMemory_155 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  DMemory_156 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  DMemory_157 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  DMemory_158 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  DMemory_159 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  DMemory_160 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  DMemory_161 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  DMemory_162 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  DMemory_163 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  DMemory_164 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  DMemory_165 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  DMemory_166 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  DMemory_167 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  DMemory_168 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  DMemory_169 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  DMemory_170 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  DMemory_171 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  DMemory_172 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  DMemory_173 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  DMemory_174 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  DMemory_175 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  DMemory_176 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  DMemory_177 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  DMemory_178 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  DMemory_179 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  DMemory_180 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  DMemory_181 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  DMemory_182 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  DMemory_183 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  DMemory_184 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  DMemory_185 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  DMemory_186 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  DMemory_187 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  DMemory_188 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  DMemory_189 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  DMemory_190 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  DMemory_191 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  DMemory_192 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  DMemory_193 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  DMemory_194 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  DMemory_195 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  DMemory_196 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  DMemory_197 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  DMemory_198 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  DMemory_199 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  DMemory_200 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  DMemory_201 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  DMemory_202 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  DMemory_203 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  DMemory_204 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  DMemory_205 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  DMemory_206 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  DMemory_207 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  DMemory_208 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  DMemory_209 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  DMemory_210 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  DMemory_211 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  DMemory_212 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  DMemory_213 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  DMemory_214 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  DMemory_215 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  DMemory_216 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  DMemory_217 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  DMemory_218 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  DMemory_219 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  DMemory_220 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  DMemory_221 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  DMemory_222 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  DMemory_223 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  DMemory_224 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  DMemory_225 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  DMemory_226 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  DMemory_227 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  DMemory_228 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  DMemory_229 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  DMemory_230 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  DMemory_231 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  DMemory_232 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  DMemory_233 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  DMemory_234 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  DMemory_235 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  DMemory_236 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  DMemory_237 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  DMemory_238 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  DMemory_239 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  DMemory_240 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  DMemory_241 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  DMemory_242 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  DMemory_243 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  DMemory_244 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  DMemory_245 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  DMemory_246 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  DMemory_247 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  DMemory_248 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  DMemory_249 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  DMemory_250 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  DMemory_251 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  DMemory_252 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  DMemory_253 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  DMemory_254 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  DMemory_255 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  DMemory_256 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  DMemory_257 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  DMemory_258 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  DMemory_259 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  DMemory_260 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  DMemory_261 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  DMemory_262 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  DMemory_263 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  DMemory_264 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  DMemory_265 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  DMemory_266 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  DMemory_267 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  DMemory_268 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  DMemory_269 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  DMemory_270 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  DMemory_271 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  DMemory_272 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  DMemory_273 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  DMemory_274 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  DMemory_275 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  DMemory_276 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  DMemory_277 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  DMemory_278 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  DMemory_279 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  DMemory_280 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  DMemory_281 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  DMemory_282 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  DMemory_283 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  DMemory_284 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  DMemory_285 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  DMemory_286 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  DMemory_287 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  DMemory_288 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  DMemory_289 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  DMemory_290 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  DMemory_291 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  DMemory_292 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  DMemory_293 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  DMemory_294 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  DMemory_295 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  DMemory_296 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  DMemory_297 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  DMemory_298 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  DMemory_299 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  DMemory_300 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  DMemory_301 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  DMemory_302 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  DMemory_303 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  DMemory_304 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  DMemory_305 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  DMemory_306 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  DMemory_307 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  DMemory_308 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  DMemory_309 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  DMemory_310 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  DMemory_311 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  DMemory_312 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  DMemory_313 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  DMemory_314 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  DMemory_315 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  DMemory_316 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  DMemory_317 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  DMemory_318 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  DMemory_319 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  DMemory_320 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  DMemory_321 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  DMemory_322 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  DMemory_323 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  DMemory_324 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  DMemory_325 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  DMemory_326 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  DMemory_327 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  DMemory_328 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  DMemory_329 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  DMemory_330 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  DMemory_331 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  DMemory_332 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  DMemory_333 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  DMemory_334 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  DMemory_335 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  DMemory_336 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  DMemory_337 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  DMemory_338 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  DMemory_339 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  DMemory_340 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  DMemory_341 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  DMemory_342 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  DMemory_343 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  DMemory_344 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  DMemory_345 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  DMemory_346 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  DMemory_347 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  DMemory_348 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  DMemory_349 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  DMemory_350 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  DMemory_351 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  DMemory_352 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  DMemory_353 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  DMemory_354 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  DMemory_355 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  DMemory_356 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  DMemory_357 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  DMemory_358 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  DMemory_359 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  DMemory_360 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  DMemory_361 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  DMemory_362 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  DMemory_363 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  DMemory_364 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  DMemory_365 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  DMemory_366 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  DMemory_367 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  DMemory_368 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  DMemory_369 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  DMemory_370 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  DMemory_371 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  DMemory_372 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  DMemory_373 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  DMemory_374 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  DMemory_375 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  DMemory_376 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  DMemory_377 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  DMemory_378 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  DMemory_379 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  DMemory_380 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  DMemory_381 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  DMemory_382 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  DMemory_383 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  DMemory_384 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  DMemory_385 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  DMemory_386 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  DMemory_387 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  DMemory_388 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  DMemory_389 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  DMemory_390 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  DMemory_391 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  DMemory_392 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  DMemory_393 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  DMemory_394 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  DMemory_395 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  DMemory_396 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  DMemory_397 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  DMemory_398 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  DMemory_399 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  DMemory_400 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  DMemory_401 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  DMemory_402 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  DMemory_403 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  DMemory_404 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  DMemory_405 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  DMemory_406 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  DMemory_407 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  DMemory_408 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  DMemory_409 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  DMemory_410 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  DMemory_411 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  DMemory_412 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  DMemory_413 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  DMemory_414 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  DMemory_415 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  DMemory_416 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  DMemory_417 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  DMemory_418 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  DMemory_419 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  DMemory_420 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  DMemory_421 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  DMemory_422 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  DMemory_423 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  DMemory_424 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  DMemory_425 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  DMemory_426 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  DMemory_427 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  DMemory_428 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  DMemory_429 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  DMemory_430 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  DMemory_431 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  DMemory_432 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  DMemory_433 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  DMemory_434 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  DMemory_435 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  DMemory_436 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  DMemory_437 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  DMemory_438 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  DMemory_439 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  DMemory_440 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  DMemory_441 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  DMemory_442 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  DMemory_443 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  DMemory_444 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  DMemory_445 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  DMemory_446 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  DMemory_447 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  DMemory_448 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  DMemory_449 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  DMemory_450 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  DMemory_451 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  DMemory_452 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  DMemory_453 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  DMemory_454 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  DMemory_455 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  DMemory_456 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  DMemory_457 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  DMemory_458 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  DMemory_459 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  DMemory_460 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  DMemory_461 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  DMemory_462 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  DMemory_463 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  DMemory_464 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  DMemory_465 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  DMemory_466 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  DMemory_467 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  DMemory_468 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  DMemory_469 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  DMemory_470 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  DMemory_471 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  DMemory_472 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  DMemory_473 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  DMemory_474 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  DMemory_475 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  DMemory_476 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  DMemory_477 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  DMemory_478 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  DMemory_479 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  DMemory_480 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  DMemory_481 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  DMemory_482 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  DMemory_483 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  DMemory_484 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  DMemory_485 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  DMemory_486 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  DMemory_487 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  DMemory_488 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  DMemory_489 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  DMemory_490 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  DMemory_491 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  DMemory_492 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  DMemory_493 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  DMemory_494 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  DMemory_495 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  DMemory_496 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  DMemory_497 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  DMemory_498 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  DMemory_499 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  DMemory_500 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  DMemory_501 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  DMemory_502 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  DMemory_503 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  DMemory_504 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  DMemory_505 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  DMemory_506 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  DMemory_507 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  DMemory_508 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  DMemory_509 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  DMemory_510 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  DMemory_511 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  DMemory_512 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  DMemory_513 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  DMemory_514 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  DMemory_515 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  DMemory_516 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  DMemory_517 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  DMemory_518 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  DMemory_519 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  DMemory_520 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  DMemory_521 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  DMemory_522 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  DMemory_523 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  DMemory_524 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  DMemory_525 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  DMemory_526 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  DMemory_527 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  DMemory_528 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  DMemory_529 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  DMemory_530 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  DMemory_531 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  DMemory_532 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  DMemory_533 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  DMemory_534 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  DMemory_535 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  DMemory_536 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  DMemory_537 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  DMemory_538 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  DMemory_539 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  DMemory_540 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  DMemory_541 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  DMemory_542 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  DMemory_543 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  DMemory_544 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  DMemory_545 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  DMemory_546 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  DMemory_547 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  DMemory_548 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  DMemory_549 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  DMemory_550 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  DMemory_551 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  DMemory_552 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  DMemory_553 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  DMemory_554 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  DMemory_555 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  DMemory_556 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  DMemory_557 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  DMemory_558 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  DMemory_559 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  DMemory_560 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  DMemory_561 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  DMemory_562 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  DMemory_563 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  DMemory_564 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  DMemory_565 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  DMemory_566 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  DMemory_567 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  DMemory_568 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  DMemory_569 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  DMemory_570 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  DMemory_571 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  DMemory_572 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  DMemory_573 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  DMemory_574 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  DMemory_575 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  DMemory_576 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  DMemory_577 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  DMemory_578 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  DMemory_579 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  DMemory_580 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  DMemory_581 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  DMemory_582 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  DMemory_583 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  DMemory_584 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  DMemory_585 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  DMemory_586 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  DMemory_587 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  DMemory_588 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  DMemory_589 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  DMemory_590 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  DMemory_591 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  DMemory_592 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  DMemory_593 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  DMemory_594 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  DMemory_595 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  DMemory_596 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  DMemory_597 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  DMemory_598 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  DMemory_599 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  DMemory_600 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  DMemory_601 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  DMemory_602 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  DMemory_603 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  DMemory_604 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  DMemory_605 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  DMemory_606 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  DMemory_607 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  DMemory_608 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  DMemory_609 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  DMemory_610 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  DMemory_611 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  DMemory_612 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  DMemory_613 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  DMemory_614 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  DMemory_615 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  DMemory_616 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  DMemory_617 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  DMemory_618 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  DMemory_619 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  DMemory_620 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  DMemory_621 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  DMemory_622 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  DMemory_623 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  DMemory_624 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  DMemory_625 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  DMemory_626 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  DMemory_627 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  DMemory_628 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  DMemory_629 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  DMemory_630 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  DMemory_631 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  DMemory_632 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  DMemory_633 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  DMemory_634 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  DMemory_635 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  DMemory_636 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  DMemory_637 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  DMemory_638 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  DMemory_639 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  DMemory_640 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  DMemory_641 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  DMemory_642 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  DMemory_643 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  DMemory_644 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  DMemory_645 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  DMemory_646 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  DMemory_647 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  DMemory_648 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  DMemory_649 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  DMemory_650 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  DMemory_651 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  DMemory_652 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  DMemory_653 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  DMemory_654 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  DMemory_655 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  DMemory_656 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  DMemory_657 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  DMemory_658 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  DMemory_659 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  DMemory_660 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  DMemory_661 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  DMemory_662 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  DMemory_663 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  DMemory_664 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  DMemory_665 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  DMemory_666 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  DMemory_667 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  DMemory_668 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  DMemory_669 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  DMemory_670 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  DMemory_671 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  DMemory_672 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  DMemory_673 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  DMemory_674 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  DMemory_675 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  DMemory_676 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  DMemory_677 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  DMemory_678 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  DMemory_679 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  DMemory_680 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  DMemory_681 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  DMemory_682 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  DMemory_683 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  DMemory_684 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  DMemory_685 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  DMemory_686 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  DMemory_687 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  DMemory_688 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  DMemory_689 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  DMemory_690 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  DMemory_691 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  DMemory_692 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  DMemory_693 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  DMemory_694 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  DMemory_695 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  DMemory_696 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  DMemory_697 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  DMemory_698 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  DMemory_699 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  DMemory_700 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  DMemory_701 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  DMemory_702 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  DMemory_703 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  DMemory_704 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  DMemory_705 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  DMemory_706 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  DMemory_707 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  DMemory_708 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  DMemory_709 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  DMemory_710 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  DMemory_711 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  DMemory_712 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  DMemory_713 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  DMemory_714 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  DMemory_715 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  DMemory_716 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  DMemory_717 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  DMemory_718 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  DMemory_719 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  DMemory_720 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  DMemory_721 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  DMemory_722 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  DMemory_723 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  DMemory_724 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  DMemory_725 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  DMemory_726 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  DMemory_727 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  DMemory_728 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  DMemory_729 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  DMemory_730 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  DMemory_731 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  DMemory_732 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  DMemory_733 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  DMemory_734 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  DMemory_735 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  DMemory_736 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  DMemory_737 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  DMemory_738 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  DMemory_739 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  DMemory_740 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  DMemory_741 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  DMemory_742 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  DMemory_743 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  DMemory_744 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  DMemory_745 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  DMemory_746 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  DMemory_747 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  DMemory_748 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  DMemory_749 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  DMemory_750 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  DMemory_751 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  DMemory_752 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  DMemory_753 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  DMemory_754 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  DMemory_755 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  DMemory_756 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  DMemory_757 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  DMemory_758 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  DMemory_759 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  DMemory_760 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  DMemory_761 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  DMemory_762 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  DMemory_763 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  DMemory_764 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  DMemory_765 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  DMemory_766 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  DMemory_767 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  DMemory_768 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  DMemory_769 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  DMemory_770 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  DMemory_771 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  DMemory_772 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  DMemory_773 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  DMemory_774 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  DMemory_775 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  DMemory_776 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  DMemory_777 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  DMemory_778 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  DMemory_779 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  DMemory_780 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  DMemory_781 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  DMemory_782 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  DMemory_783 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  DMemory_784 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  DMemory_785 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  DMemory_786 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  DMemory_787 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  DMemory_788 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  DMemory_789 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  DMemory_790 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  DMemory_791 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  DMemory_792 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  DMemory_793 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  DMemory_794 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  DMemory_795 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  DMemory_796 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  DMemory_797 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  DMemory_798 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  DMemory_799 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  DMemory_800 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  DMemory_801 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  DMemory_802 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  DMemory_803 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  DMemory_804 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  DMemory_805 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  DMemory_806 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  DMemory_807 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  DMemory_808 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  DMemory_809 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  DMemory_810 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  DMemory_811 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  DMemory_812 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  DMemory_813 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  DMemory_814 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  DMemory_815 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  DMemory_816 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  DMemory_817 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  DMemory_818 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  DMemory_819 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  DMemory_820 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  DMemory_821 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  DMemory_822 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  DMemory_823 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  DMemory_824 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  DMemory_825 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  DMemory_826 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  DMemory_827 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  DMemory_828 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  DMemory_829 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  DMemory_830 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  DMemory_831 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  DMemory_832 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  DMemory_833 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  DMemory_834 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  DMemory_835 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  DMemory_836 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  DMemory_837 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  DMemory_838 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  DMemory_839 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  DMemory_840 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  DMemory_841 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  DMemory_842 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  DMemory_843 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  DMemory_844 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  DMemory_845 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  DMemory_846 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  DMemory_847 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  DMemory_848 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  DMemory_849 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  DMemory_850 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  DMemory_851 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  DMemory_852 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  DMemory_853 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  DMemory_854 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  DMemory_855 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  DMemory_856 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  DMemory_857 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  DMemory_858 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  DMemory_859 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  DMemory_860 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  DMemory_861 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  DMemory_862 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  DMemory_863 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  DMemory_864 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  DMemory_865 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  DMemory_866 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  DMemory_867 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  DMemory_868 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  DMemory_869 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  DMemory_870 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  DMemory_871 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  DMemory_872 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  DMemory_873 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  DMemory_874 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  DMemory_875 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  DMemory_876 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  DMemory_877 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  DMemory_878 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  DMemory_879 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  DMemory_880 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  DMemory_881 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  DMemory_882 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  DMemory_883 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  DMemory_884 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  DMemory_885 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  DMemory_886 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  DMemory_887 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  DMemory_888 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  DMemory_889 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  DMemory_890 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  DMemory_891 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  DMemory_892 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  DMemory_893 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  DMemory_894 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  DMemory_895 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  DMemory_896 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  DMemory_897 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  DMemory_898 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  DMemory_899 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  DMemory_900 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  DMemory_901 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  DMemory_902 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  DMemory_903 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  DMemory_904 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  DMemory_905 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  DMemory_906 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  DMemory_907 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  DMemory_908 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  DMemory_909 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  DMemory_910 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  DMemory_911 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  DMemory_912 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  DMemory_913 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  DMemory_914 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  DMemory_915 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  DMemory_916 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  DMemory_917 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  DMemory_918 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  DMemory_919 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  DMemory_920 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  DMemory_921 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  DMemory_922 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  DMemory_923 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  DMemory_924 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  DMemory_925 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  DMemory_926 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  DMemory_927 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  DMemory_928 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  DMemory_929 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  DMemory_930 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  DMemory_931 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  DMemory_932 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  DMemory_933 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  DMemory_934 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  DMemory_935 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  DMemory_936 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  DMemory_937 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  DMemory_938 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  DMemory_939 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  DMemory_940 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  DMemory_941 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  DMemory_942 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  DMemory_943 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  DMemory_944 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  DMemory_945 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  DMemory_946 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  DMemory_947 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  DMemory_948 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  DMemory_949 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  DMemory_950 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  DMemory_951 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  DMemory_952 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  DMemory_953 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  DMemory_954 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  DMemory_955 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  DMemory_956 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  DMemory_957 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  DMemory_958 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  DMemory_959 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  DMemory_960 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  DMemory_961 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  DMemory_962 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  DMemory_963 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  DMemory_964 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  DMemory_965 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  DMemory_966 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  DMemory_967 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  DMemory_968 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  DMemory_969 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  DMemory_970 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  DMemory_971 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  DMemory_972 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  DMemory_973 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  DMemory_974 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  DMemory_975 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  DMemory_976 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  DMemory_977 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  DMemory_978 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  DMemory_979 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  DMemory_980 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  DMemory_981 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  DMemory_982 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  DMemory_983 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  DMemory_984 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  DMemory_985 = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  DMemory_986 = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  DMemory_987 = _RAND_1025[31:0];
  _RAND_1026 = {1{`RANDOM}};
  DMemory_988 = _RAND_1026[31:0];
  _RAND_1027 = {1{`RANDOM}};
  DMemory_989 = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  DMemory_990 = _RAND_1028[31:0];
  _RAND_1029 = {1{`RANDOM}};
  DMemory_991 = _RAND_1029[31:0];
  _RAND_1030 = {1{`RANDOM}};
  DMemory_992 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  DMemory_993 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  DMemory_994 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  DMemory_995 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  DMemory_996 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  DMemory_997 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  DMemory_998 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  DMemory_999 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  DMemory_1000 = _RAND_1038[31:0];
  _RAND_1039 = {1{`RANDOM}};
  DMemory_1001 = _RAND_1039[31:0];
  _RAND_1040 = {1{`RANDOM}};
  DMemory_1002 = _RAND_1040[31:0];
  _RAND_1041 = {1{`RANDOM}};
  DMemory_1003 = _RAND_1041[31:0];
  _RAND_1042 = {1{`RANDOM}};
  DMemory_1004 = _RAND_1042[31:0];
  _RAND_1043 = {1{`RANDOM}};
  DMemory_1005 = _RAND_1043[31:0];
  _RAND_1044 = {1{`RANDOM}};
  DMemory_1006 = _RAND_1044[31:0];
  _RAND_1045 = {1{`RANDOM}};
  DMemory_1007 = _RAND_1045[31:0];
  _RAND_1046 = {1{`RANDOM}};
  DMemory_1008 = _RAND_1046[31:0];
  _RAND_1047 = {1{`RANDOM}};
  DMemory_1009 = _RAND_1047[31:0];
  _RAND_1048 = {1{`RANDOM}};
  DMemory_1010 = _RAND_1048[31:0];
  _RAND_1049 = {1{`RANDOM}};
  DMemory_1011 = _RAND_1049[31:0];
  _RAND_1050 = {1{`RANDOM}};
  DMemory_1012 = _RAND_1050[31:0];
  _RAND_1051 = {1{`RANDOM}};
  DMemory_1013 = _RAND_1051[31:0];
  _RAND_1052 = {1{`RANDOM}};
  DMemory_1014 = _RAND_1052[31:0];
  _RAND_1053 = {1{`RANDOM}};
  DMemory_1015 = _RAND_1053[31:0];
  _RAND_1054 = {1{`RANDOM}};
  DMemory_1016 = _RAND_1054[31:0];
  _RAND_1055 = {1{`RANDOM}};
  DMemory_1017 = _RAND_1055[31:0];
  _RAND_1056 = {1{`RANDOM}};
  DMemory_1018 = _RAND_1056[31:0];
  _RAND_1057 = {1{`RANDOM}};
  DMemory_1019 = _RAND_1057[31:0];
  _RAND_1058 = {1{`RANDOM}};
  DMemory_1020 = _RAND_1058[31:0];
  _RAND_1059 = {1{`RANDOM}};
  DMemory_1021 = _RAND_1059[31:0];
  _RAND_1060 = {1{`RANDOM}};
  DMemory_1022 = _RAND_1060[31:0];
  _RAND_1061 = {1{`RANDOM}};
  DMemory_1023 = _RAND_1061[31:0];
  _RAND_1062 = {1{`RANDOM}};
  IMemory_0 = _RAND_1062[31:0];
  _RAND_1063 = {1{`RANDOM}};
  IMemory_1 = _RAND_1063[31:0];
  _RAND_1064 = {1{`RANDOM}};
  IFIDIR = _RAND_1064[31:0];
  _RAND_1065 = {1{`RANDOM}};
  IDEXIR = _RAND_1065[31:0];
  _RAND_1066 = {1{`RANDOM}};
  EXMEMIR = _RAND_1066[31:0];
  _RAND_1067 = {1{`RANDOM}};
  MEMWBIR = _RAND_1067[31:0];
  _RAND_1068 = {2{`RANDOM}};
  CurPC = _RAND_1068[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ControlUnit(
  input         clock,
  input         reset,
  input         io_reset,
  input  [31:0] io_insns_0,
  input  [31:0] io_insns_1,
  input  [63:0] io_PC,
  output [63:0] io_nPC,
  output [31:0] io_insn
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] counterReg; // @[cpu.scala 37:27]
  wire [1:0] _counterReg_T_1 = counterReg + 2'h1; // @[cpu.scala 41:30]
  wire [63:0] _io_nPC_T_1 = io_PC + 64'h4; // @[cpu.scala 44:21]
  wire [63:0] _io_insn_T = {{2'd0}, io_PC[63:2]}; // @[cpu.scala 45:32]
  wire [31:0] _GEN_2 = 10'h1 == _io_insn_T[9:0] ? io_insns_1 : io_insns_0; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_3 = 10'h2 == _io_insn_T[9:0] ? 32'h13 : _GEN_2; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_4 = 10'h3 == _io_insn_T[9:0] ? 32'h13 : _GEN_3; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_5 = 10'h4 == _io_insn_T[9:0] ? 32'h13 : _GEN_4; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_6 = 10'h5 == _io_insn_T[9:0] ? 32'h13 : _GEN_5; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_7 = 10'h6 == _io_insn_T[9:0] ? 32'h13 : _GEN_6; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_8 = 10'h7 == _io_insn_T[9:0] ? 32'h13 : _GEN_7; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_9 = 10'h8 == _io_insn_T[9:0] ? 32'h13 : _GEN_8; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_10 = 10'h9 == _io_insn_T[9:0] ? 32'h13 : _GEN_9; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_11 = 10'ha == _io_insn_T[9:0] ? 32'h13 : _GEN_10; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_12 = 10'hb == _io_insn_T[9:0] ? 32'h13 : _GEN_11; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_13 = 10'hc == _io_insn_T[9:0] ? 32'h13 : _GEN_12; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_14 = 10'hd == _io_insn_T[9:0] ? 32'h13 : _GEN_13; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_15 = 10'he == _io_insn_T[9:0] ? 32'h13 : _GEN_14; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_16 = 10'hf == _io_insn_T[9:0] ? 32'h13 : _GEN_15; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_17 = 10'h10 == _io_insn_T[9:0] ? 32'h13 : _GEN_16; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_18 = 10'h11 == _io_insn_T[9:0] ? 32'h13 : _GEN_17; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_19 = 10'h12 == _io_insn_T[9:0] ? 32'h13 : _GEN_18; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_20 = 10'h13 == _io_insn_T[9:0] ? 32'h13 : _GEN_19; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_21 = 10'h14 == _io_insn_T[9:0] ? 32'h13 : _GEN_20; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_22 = 10'h15 == _io_insn_T[9:0] ? 32'h13 : _GEN_21; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_23 = 10'h16 == _io_insn_T[9:0] ? 32'h13 : _GEN_22; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_24 = 10'h17 == _io_insn_T[9:0] ? 32'h13 : _GEN_23; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_25 = 10'h18 == _io_insn_T[9:0] ? 32'h13 : _GEN_24; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_26 = 10'h19 == _io_insn_T[9:0] ? 32'h13 : _GEN_25; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_27 = 10'h1a == _io_insn_T[9:0] ? 32'h13 : _GEN_26; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_28 = 10'h1b == _io_insn_T[9:0] ? 32'h13 : _GEN_27; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_29 = 10'h1c == _io_insn_T[9:0] ? 32'h13 : _GEN_28; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_30 = 10'h1d == _io_insn_T[9:0] ? 32'h13 : _GEN_29; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_31 = 10'h1e == _io_insn_T[9:0] ? 32'h13 : _GEN_30; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_32 = 10'h1f == _io_insn_T[9:0] ? 32'h13 : _GEN_31; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_33 = 10'h20 == _io_insn_T[9:0] ? 32'h13 : _GEN_32; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_34 = 10'h21 == _io_insn_T[9:0] ? 32'h13 : _GEN_33; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_35 = 10'h22 == _io_insn_T[9:0] ? 32'h13 : _GEN_34; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_36 = 10'h23 == _io_insn_T[9:0] ? 32'h13 : _GEN_35; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_37 = 10'h24 == _io_insn_T[9:0] ? 32'h13 : _GEN_36; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_38 = 10'h25 == _io_insn_T[9:0] ? 32'h13 : _GEN_37; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_39 = 10'h26 == _io_insn_T[9:0] ? 32'h13 : _GEN_38; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_40 = 10'h27 == _io_insn_T[9:0] ? 32'h13 : _GEN_39; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_41 = 10'h28 == _io_insn_T[9:0] ? 32'h13 : _GEN_40; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_42 = 10'h29 == _io_insn_T[9:0] ? 32'h13 : _GEN_41; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_43 = 10'h2a == _io_insn_T[9:0] ? 32'h13 : _GEN_42; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_44 = 10'h2b == _io_insn_T[9:0] ? 32'h13 : _GEN_43; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_45 = 10'h2c == _io_insn_T[9:0] ? 32'h13 : _GEN_44; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_46 = 10'h2d == _io_insn_T[9:0] ? 32'h13 : _GEN_45; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_47 = 10'h2e == _io_insn_T[9:0] ? 32'h13 : _GEN_46; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_48 = 10'h2f == _io_insn_T[9:0] ? 32'h13 : _GEN_47; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_49 = 10'h30 == _io_insn_T[9:0] ? 32'h13 : _GEN_48; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_50 = 10'h31 == _io_insn_T[9:0] ? 32'h13 : _GEN_49; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_51 = 10'h32 == _io_insn_T[9:0] ? 32'h13 : _GEN_50; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_52 = 10'h33 == _io_insn_T[9:0] ? 32'h13 : _GEN_51; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_53 = 10'h34 == _io_insn_T[9:0] ? 32'h13 : _GEN_52; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_54 = 10'h35 == _io_insn_T[9:0] ? 32'h13 : _GEN_53; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_55 = 10'h36 == _io_insn_T[9:0] ? 32'h13 : _GEN_54; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_56 = 10'h37 == _io_insn_T[9:0] ? 32'h13 : _GEN_55; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_57 = 10'h38 == _io_insn_T[9:0] ? 32'h13 : _GEN_56; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_58 = 10'h39 == _io_insn_T[9:0] ? 32'h13 : _GEN_57; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_59 = 10'h3a == _io_insn_T[9:0] ? 32'h13 : _GEN_58; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_60 = 10'h3b == _io_insn_T[9:0] ? 32'h13 : _GEN_59; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_61 = 10'h3c == _io_insn_T[9:0] ? 32'h13 : _GEN_60; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_62 = 10'h3d == _io_insn_T[9:0] ? 32'h13 : _GEN_61; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_63 = 10'h3e == _io_insn_T[9:0] ? 32'h13 : _GEN_62; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_64 = 10'h3f == _io_insn_T[9:0] ? 32'h13 : _GEN_63; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_65 = 10'h40 == _io_insn_T[9:0] ? 32'h13 : _GEN_64; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_66 = 10'h41 == _io_insn_T[9:0] ? 32'h13 : _GEN_65; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_67 = 10'h42 == _io_insn_T[9:0] ? 32'h13 : _GEN_66; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_68 = 10'h43 == _io_insn_T[9:0] ? 32'h13 : _GEN_67; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_69 = 10'h44 == _io_insn_T[9:0] ? 32'h13 : _GEN_68; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_70 = 10'h45 == _io_insn_T[9:0] ? 32'h13 : _GEN_69; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_71 = 10'h46 == _io_insn_T[9:0] ? 32'h13 : _GEN_70; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_72 = 10'h47 == _io_insn_T[9:0] ? 32'h13 : _GEN_71; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_73 = 10'h48 == _io_insn_T[9:0] ? 32'h13 : _GEN_72; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_74 = 10'h49 == _io_insn_T[9:0] ? 32'h13 : _GEN_73; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_75 = 10'h4a == _io_insn_T[9:0] ? 32'h13 : _GEN_74; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_76 = 10'h4b == _io_insn_T[9:0] ? 32'h13 : _GEN_75; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_77 = 10'h4c == _io_insn_T[9:0] ? 32'h13 : _GEN_76; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_78 = 10'h4d == _io_insn_T[9:0] ? 32'h13 : _GEN_77; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_79 = 10'h4e == _io_insn_T[9:0] ? 32'h13 : _GEN_78; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_80 = 10'h4f == _io_insn_T[9:0] ? 32'h13 : _GEN_79; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_81 = 10'h50 == _io_insn_T[9:0] ? 32'h13 : _GEN_80; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_82 = 10'h51 == _io_insn_T[9:0] ? 32'h13 : _GEN_81; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_83 = 10'h52 == _io_insn_T[9:0] ? 32'h13 : _GEN_82; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_84 = 10'h53 == _io_insn_T[9:0] ? 32'h13 : _GEN_83; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_85 = 10'h54 == _io_insn_T[9:0] ? 32'h13 : _GEN_84; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_86 = 10'h55 == _io_insn_T[9:0] ? 32'h13 : _GEN_85; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_87 = 10'h56 == _io_insn_T[9:0] ? 32'h13 : _GEN_86; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_88 = 10'h57 == _io_insn_T[9:0] ? 32'h13 : _GEN_87; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_89 = 10'h58 == _io_insn_T[9:0] ? 32'h13 : _GEN_88; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_90 = 10'h59 == _io_insn_T[9:0] ? 32'h13 : _GEN_89; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_91 = 10'h5a == _io_insn_T[9:0] ? 32'h13 : _GEN_90; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_92 = 10'h5b == _io_insn_T[9:0] ? 32'h13 : _GEN_91; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_93 = 10'h5c == _io_insn_T[9:0] ? 32'h13 : _GEN_92; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_94 = 10'h5d == _io_insn_T[9:0] ? 32'h13 : _GEN_93; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_95 = 10'h5e == _io_insn_T[9:0] ? 32'h13 : _GEN_94; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_96 = 10'h5f == _io_insn_T[9:0] ? 32'h13 : _GEN_95; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_97 = 10'h60 == _io_insn_T[9:0] ? 32'h13 : _GEN_96; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_98 = 10'h61 == _io_insn_T[9:0] ? 32'h13 : _GEN_97; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_99 = 10'h62 == _io_insn_T[9:0] ? 32'h13 : _GEN_98; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_100 = 10'h63 == _io_insn_T[9:0] ? 32'h13 : _GEN_99; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_101 = 10'h64 == _io_insn_T[9:0] ? 32'h13 : _GEN_100; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_102 = 10'h65 == _io_insn_T[9:0] ? 32'h13 : _GEN_101; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_103 = 10'h66 == _io_insn_T[9:0] ? 32'h13 : _GEN_102; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_104 = 10'h67 == _io_insn_T[9:0] ? 32'h13 : _GEN_103; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_105 = 10'h68 == _io_insn_T[9:0] ? 32'h13 : _GEN_104; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_106 = 10'h69 == _io_insn_T[9:0] ? 32'h13 : _GEN_105; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_107 = 10'h6a == _io_insn_T[9:0] ? 32'h13 : _GEN_106; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_108 = 10'h6b == _io_insn_T[9:0] ? 32'h13 : _GEN_107; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_109 = 10'h6c == _io_insn_T[9:0] ? 32'h13 : _GEN_108; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_110 = 10'h6d == _io_insn_T[9:0] ? 32'h13 : _GEN_109; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_111 = 10'h6e == _io_insn_T[9:0] ? 32'h13 : _GEN_110; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_112 = 10'h6f == _io_insn_T[9:0] ? 32'h13 : _GEN_111; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_113 = 10'h70 == _io_insn_T[9:0] ? 32'h13 : _GEN_112; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_114 = 10'h71 == _io_insn_T[9:0] ? 32'h13 : _GEN_113; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_115 = 10'h72 == _io_insn_T[9:0] ? 32'h13 : _GEN_114; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_116 = 10'h73 == _io_insn_T[9:0] ? 32'h13 : _GEN_115; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_117 = 10'h74 == _io_insn_T[9:0] ? 32'h13 : _GEN_116; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_118 = 10'h75 == _io_insn_T[9:0] ? 32'h13 : _GEN_117; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_119 = 10'h76 == _io_insn_T[9:0] ? 32'h13 : _GEN_118; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_120 = 10'h77 == _io_insn_T[9:0] ? 32'h13 : _GEN_119; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_121 = 10'h78 == _io_insn_T[9:0] ? 32'h13 : _GEN_120; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_122 = 10'h79 == _io_insn_T[9:0] ? 32'h13 : _GEN_121; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_123 = 10'h7a == _io_insn_T[9:0] ? 32'h13 : _GEN_122; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_124 = 10'h7b == _io_insn_T[9:0] ? 32'h13 : _GEN_123; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_125 = 10'h7c == _io_insn_T[9:0] ? 32'h13 : _GEN_124; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_126 = 10'h7d == _io_insn_T[9:0] ? 32'h13 : _GEN_125; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_127 = 10'h7e == _io_insn_T[9:0] ? 32'h13 : _GEN_126; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_128 = 10'h7f == _io_insn_T[9:0] ? 32'h13 : _GEN_127; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_129 = 10'h80 == _io_insn_T[9:0] ? 32'h13 : _GEN_128; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_130 = 10'h81 == _io_insn_T[9:0] ? 32'h13 : _GEN_129; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_131 = 10'h82 == _io_insn_T[9:0] ? 32'h13 : _GEN_130; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_132 = 10'h83 == _io_insn_T[9:0] ? 32'h13 : _GEN_131; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_133 = 10'h84 == _io_insn_T[9:0] ? 32'h13 : _GEN_132; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_134 = 10'h85 == _io_insn_T[9:0] ? 32'h13 : _GEN_133; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_135 = 10'h86 == _io_insn_T[9:0] ? 32'h13 : _GEN_134; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_136 = 10'h87 == _io_insn_T[9:0] ? 32'h13 : _GEN_135; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_137 = 10'h88 == _io_insn_T[9:0] ? 32'h13 : _GEN_136; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_138 = 10'h89 == _io_insn_T[9:0] ? 32'h13 : _GEN_137; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_139 = 10'h8a == _io_insn_T[9:0] ? 32'h13 : _GEN_138; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_140 = 10'h8b == _io_insn_T[9:0] ? 32'h13 : _GEN_139; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_141 = 10'h8c == _io_insn_T[9:0] ? 32'h13 : _GEN_140; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_142 = 10'h8d == _io_insn_T[9:0] ? 32'h13 : _GEN_141; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_143 = 10'h8e == _io_insn_T[9:0] ? 32'h13 : _GEN_142; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_144 = 10'h8f == _io_insn_T[9:0] ? 32'h13 : _GEN_143; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_145 = 10'h90 == _io_insn_T[9:0] ? 32'h13 : _GEN_144; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_146 = 10'h91 == _io_insn_T[9:0] ? 32'h13 : _GEN_145; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_147 = 10'h92 == _io_insn_T[9:0] ? 32'h13 : _GEN_146; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_148 = 10'h93 == _io_insn_T[9:0] ? 32'h13 : _GEN_147; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_149 = 10'h94 == _io_insn_T[9:0] ? 32'h13 : _GEN_148; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_150 = 10'h95 == _io_insn_T[9:0] ? 32'h13 : _GEN_149; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_151 = 10'h96 == _io_insn_T[9:0] ? 32'h13 : _GEN_150; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_152 = 10'h97 == _io_insn_T[9:0] ? 32'h13 : _GEN_151; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_153 = 10'h98 == _io_insn_T[9:0] ? 32'h13 : _GEN_152; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_154 = 10'h99 == _io_insn_T[9:0] ? 32'h13 : _GEN_153; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_155 = 10'h9a == _io_insn_T[9:0] ? 32'h13 : _GEN_154; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_156 = 10'h9b == _io_insn_T[9:0] ? 32'h13 : _GEN_155; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_157 = 10'h9c == _io_insn_T[9:0] ? 32'h13 : _GEN_156; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_158 = 10'h9d == _io_insn_T[9:0] ? 32'h13 : _GEN_157; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_159 = 10'h9e == _io_insn_T[9:0] ? 32'h13 : _GEN_158; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_160 = 10'h9f == _io_insn_T[9:0] ? 32'h13 : _GEN_159; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_161 = 10'ha0 == _io_insn_T[9:0] ? 32'h13 : _GEN_160; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_162 = 10'ha1 == _io_insn_T[9:0] ? 32'h13 : _GEN_161; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_163 = 10'ha2 == _io_insn_T[9:0] ? 32'h13 : _GEN_162; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_164 = 10'ha3 == _io_insn_T[9:0] ? 32'h13 : _GEN_163; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_165 = 10'ha4 == _io_insn_T[9:0] ? 32'h13 : _GEN_164; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_166 = 10'ha5 == _io_insn_T[9:0] ? 32'h13 : _GEN_165; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_167 = 10'ha6 == _io_insn_T[9:0] ? 32'h13 : _GEN_166; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_168 = 10'ha7 == _io_insn_T[9:0] ? 32'h13 : _GEN_167; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_169 = 10'ha8 == _io_insn_T[9:0] ? 32'h13 : _GEN_168; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_170 = 10'ha9 == _io_insn_T[9:0] ? 32'h13 : _GEN_169; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_171 = 10'haa == _io_insn_T[9:0] ? 32'h13 : _GEN_170; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_172 = 10'hab == _io_insn_T[9:0] ? 32'h13 : _GEN_171; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_173 = 10'hac == _io_insn_T[9:0] ? 32'h13 : _GEN_172; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_174 = 10'had == _io_insn_T[9:0] ? 32'h13 : _GEN_173; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_175 = 10'hae == _io_insn_T[9:0] ? 32'h13 : _GEN_174; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_176 = 10'haf == _io_insn_T[9:0] ? 32'h13 : _GEN_175; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_177 = 10'hb0 == _io_insn_T[9:0] ? 32'h13 : _GEN_176; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_178 = 10'hb1 == _io_insn_T[9:0] ? 32'h13 : _GEN_177; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_179 = 10'hb2 == _io_insn_T[9:0] ? 32'h13 : _GEN_178; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_180 = 10'hb3 == _io_insn_T[9:0] ? 32'h13 : _GEN_179; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_181 = 10'hb4 == _io_insn_T[9:0] ? 32'h13 : _GEN_180; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_182 = 10'hb5 == _io_insn_T[9:0] ? 32'h13 : _GEN_181; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_183 = 10'hb6 == _io_insn_T[9:0] ? 32'h13 : _GEN_182; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_184 = 10'hb7 == _io_insn_T[9:0] ? 32'h13 : _GEN_183; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_185 = 10'hb8 == _io_insn_T[9:0] ? 32'h13 : _GEN_184; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_186 = 10'hb9 == _io_insn_T[9:0] ? 32'h13 : _GEN_185; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_187 = 10'hba == _io_insn_T[9:0] ? 32'h13 : _GEN_186; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_188 = 10'hbb == _io_insn_T[9:0] ? 32'h13 : _GEN_187; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_189 = 10'hbc == _io_insn_T[9:0] ? 32'h13 : _GEN_188; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_190 = 10'hbd == _io_insn_T[9:0] ? 32'h13 : _GEN_189; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_191 = 10'hbe == _io_insn_T[9:0] ? 32'h13 : _GEN_190; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_192 = 10'hbf == _io_insn_T[9:0] ? 32'h13 : _GEN_191; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_193 = 10'hc0 == _io_insn_T[9:0] ? 32'h13 : _GEN_192; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_194 = 10'hc1 == _io_insn_T[9:0] ? 32'h13 : _GEN_193; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_195 = 10'hc2 == _io_insn_T[9:0] ? 32'h13 : _GEN_194; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_196 = 10'hc3 == _io_insn_T[9:0] ? 32'h13 : _GEN_195; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_197 = 10'hc4 == _io_insn_T[9:0] ? 32'h13 : _GEN_196; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_198 = 10'hc5 == _io_insn_T[9:0] ? 32'h13 : _GEN_197; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_199 = 10'hc6 == _io_insn_T[9:0] ? 32'h13 : _GEN_198; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_200 = 10'hc7 == _io_insn_T[9:0] ? 32'h13 : _GEN_199; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_201 = 10'hc8 == _io_insn_T[9:0] ? 32'h13 : _GEN_200; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_202 = 10'hc9 == _io_insn_T[9:0] ? 32'h13 : _GEN_201; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_203 = 10'hca == _io_insn_T[9:0] ? 32'h13 : _GEN_202; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_204 = 10'hcb == _io_insn_T[9:0] ? 32'h13 : _GEN_203; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_205 = 10'hcc == _io_insn_T[9:0] ? 32'h13 : _GEN_204; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_206 = 10'hcd == _io_insn_T[9:0] ? 32'h13 : _GEN_205; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_207 = 10'hce == _io_insn_T[9:0] ? 32'h13 : _GEN_206; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_208 = 10'hcf == _io_insn_T[9:0] ? 32'h13 : _GEN_207; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_209 = 10'hd0 == _io_insn_T[9:0] ? 32'h13 : _GEN_208; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_210 = 10'hd1 == _io_insn_T[9:0] ? 32'h13 : _GEN_209; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_211 = 10'hd2 == _io_insn_T[9:0] ? 32'h13 : _GEN_210; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_212 = 10'hd3 == _io_insn_T[9:0] ? 32'h13 : _GEN_211; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_213 = 10'hd4 == _io_insn_T[9:0] ? 32'h13 : _GEN_212; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_214 = 10'hd5 == _io_insn_T[9:0] ? 32'h13 : _GEN_213; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_215 = 10'hd6 == _io_insn_T[9:0] ? 32'h13 : _GEN_214; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_216 = 10'hd7 == _io_insn_T[9:0] ? 32'h13 : _GEN_215; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_217 = 10'hd8 == _io_insn_T[9:0] ? 32'h13 : _GEN_216; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_218 = 10'hd9 == _io_insn_T[9:0] ? 32'h13 : _GEN_217; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_219 = 10'hda == _io_insn_T[9:0] ? 32'h13 : _GEN_218; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_220 = 10'hdb == _io_insn_T[9:0] ? 32'h13 : _GEN_219; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_221 = 10'hdc == _io_insn_T[9:0] ? 32'h13 : _GEN_220; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_222 = 10'hdd == _io_insn_T[9:0] ? 32'h13 : _GEN_221; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_223 = 10'hde == _io_insn_T[9:0] ? 32'h13 : _GEN_222; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_224 = 10'hdf == _io_insn_T[9:0] ? 32'h13 : _GEN_223; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_225 = 10'he0 == _io_insn_T[9:0] ? 32'h13 : _GEN_224; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_226 = 10'he1 == _io_insn_T[9:0] ? 32'h13 : _GEN_225; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_227 = 10'he2 == _io_insn_T[9:0] ? 32'h13 : _GEN_226; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_228 = 10'he3 == _io_insn_T[9:0] ? 32'h13 : _GEN_227; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_229 = 10'he4 == _io_insn_T[9:0] ? 32'h13 : _GEN_228; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_230 = 10'he5 == _io_insn_T[9:0] ? 32'h13 : _GEN_229; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_231 = 10'he6 == _io_insn_T[9:0] ? 32'h13 : _GEN_230; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_232 = 10'he7 == _io_insn_T[9:0] ? 32'h13 : _GEN_231; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_233 = 10'he8 == _io_insn_T[9:0] ? 32'h13 : _GEN_232; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_234 = 10'he9 == _io_insn_T[9:0] ? 32'h13 : _GEN_233; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_235 = 10'hea == _io_insn_T[9:0] ? 32'h13 : _GEN_234; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_236 = 10'heb == _io_insn_T[9:0] ? 32'h13 : _GEN_235; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_237 = 10'hec == _io_insn_T[9:0] ? 32'h13 : _GEN_236; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_238 = 10'hed == _io_insn_T[9:0] ? 32'h13 : _GEN_237; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_239 = 10'hee == _io_insn_T[9:0] ? 32'h13 : _GEN_238; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_240 = 10'hef == _io_insn_T[9:0] ? 32'h13 : _GEN_239; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_241 = 10'hf0 == _io_insn_T[9:0] ? 32'h13 : _GEN_240; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_242 = 10'hf1 == _io_insn_T[9:0] ? 32'h13 : _GEN_241; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_243 = 10'hf2 == _io_insn_T[9:0] ? 32'h13 : _GEN_242; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_244 = 10'hf3 == _io_insn_T[9:0] ? 32'h13 : _GEN_243; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_245 = 10'hf4 == _io_insn_T[9:0] ? 32'h13 : _GEN_244; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_246 = 10'hf5 == _io_insn_T[9:0] ? 32'h13 : _GEN_245; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_247 = 10'hf6 == _io_insn_T[9:0] ? 32'h13 : _GEN_246; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_248 = 10'hf7 == _io_insn_T[9:0] ? 32'h13 : _GEN_247; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_249 = 10'hf8 == _io_insn_T[9:0] ? 32'h13 : _GEN_248; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_250 = 10'hf9 == _io_insn_T[9:0] ? 32'h13 : _GEN_249; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_251 = 10'hfa == _io_insn_T[9:0] ? 32'h13 : _GEN_250; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_252 = 10'hfb == _io_insn_T[9:0] ? 32'h13 : _GEN_251; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_253 = 10'hfc == _io_insn_T[9:0] ? 32'h13 : _GEN_252; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_254 = 10'hfd == _io_insn_T[9:0] ? 32'h13 : _GEN_253; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_255 = 10'hfe == _io_insn_T[9:0] ? 32'h13 : _GEN_254; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_256 = 10'hff == _io_insn_T[9:0] ? 32'h13 : _GEN_255; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_257 = 10'h100 == _io_insn_T[9:0] ? 32'h13 : _GEN_256; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_258 = 10'h101 == _io_insn_T[9:0] ? 32'h13 : _GEN_257; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_259 = 10'h102 == _io_insn_T[9:0] ? 32'h13 : _GEN_258; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_260 = 10'h103 == _io_insn_T[9:0] ? 32'h13 : _GEN_259; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_261 = 10'h104 == _io_insn_T[9:0] ? 32'h13 : _GEN_260; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_262 = 10'h105 == _io_insn_T[9:0] ? 32'h13 : _GEN_261; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_263 = 10'h106 == _io_insn_T[9:0] ? 32'h13 : _GEN_262; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_264 = 10'h107 == _io_insn_T[9:0] ? 32'h13 : _GEN_263; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_265 = 10'h108 == _io_insn_T[9:0] ? 32'h13 : _GEN_264; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_266 = 10'h109 == _io_insn_T[9:0] ? 32'h13 : _GEN_265; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_267 = 10'h10a == _io_insn_T[9:0] ? 32'h13 : _GEN_266; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_268 = 10'h10b == _io_insn_T[9:0] ? 32'h13 : _GEN_267; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_269 = 10'h10c == _io_insn_T[9:0] ? 32'h13 : _GEN_268; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_270 = 10'h10d == _io_insn_T[9:0] ? 32'h13 : _GEN_269; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_271 = 10'h10e == _io_insn_T[9:0] ? 32'h13 : _GEN_270; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_272 = 10'h10f == _io_insn_T[9:0] ? 32'h13 : _GEN_271; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_273 = 10'h110 == _io_insn_T[9:0] ? 32'h13 : _GEN_272; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_274 = 10'h111 == _io_insn_T[9:0] ? 32'h13 : _GEN_273; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_275 = 10'h112 == _io_insn_T[9:0] ? 32'h13 : _GEN_274; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_276 = 10'h113 == _io_insn_T[9:0] ? 32'h13 : _GEN_275; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_277 = 10'h114 == _io_insn_T[9:0] ? 32'h13 : _GEN_276; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_278 = 10'h115 == _io_insn_T[9:0] ? 32'h13 : _GEN_277; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_279 = 10'h116 == _io_insn_T[9:0] ? 32'h13 : _GEN_278; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_280 = 10'h117 == _io_insn_T[9:0] ? 32'h13 : _GEN_279; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_281 = 10'h118 == _io_insn_T[9:0] ? 32'h13 : _GEN_280; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_282 = 10'h119 == _io_insn_T[9:0] ? 32'h13 : _GEN_281; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_283 = 10'h11a == _io_insn_T[9:0] ? 32'h13 : _GEN_282; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_284 = 10'h11b == _io_insn_T[9:0] ? 32'h13 : _GEN_283; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_285 = 10'h11c == _io_insn_T[9:0] ? 32'h13 : _GEN_284; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_286 = 10'h11d == _io_insn_T[9:0] ? 32'h13 : _GEN_285; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_287 = 10'h11e == _io_insn_T[9:0] ? 32'h13 : _GEN_286; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_288 = 10'h11f == _io_insn_T[9:0] ? 32'h13 : _GEN_287; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_289 = 10'h120 == _io_insn_T[9:0] ? 32'h13 : _GEN_288; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_290 = 10'h121 == _io_insn_T[9:0] ? 32'h13 : _GEN_289; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_291 = 10'h122 == _io_insn_T[9:0] ? 32'h13 : _GEN_290; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_292 = 10'h123 == _io_insn_T[9:0] ? 32'h13 : _GEN_291; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_293 = 10'h124 == _io_insn_T[9:0] ? 32'h13 : _GEN_292; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_294 = 10'h125 == _io_insn_T[9:0] ? 32'h13 : _GEN_293; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_295 = 10'h126 == _io_insn_T[9:0] ? 32'h13 : _GEN_294; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_296 = 10'h127 == _io_insn_T[9:0] ? 32'h13 : _GEN_295; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_297 = 10'h128 == _io_insn_T[9:0] ? 32'h13 : _GEN_296; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_298 = 10'h129 == _io_insn_T[9:0] ? 32'h13 : _GEN_297; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_299 = 10'h12a == _io_insn_T[9:0] ? 32'h13 : _GEN_298; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_300 = 10'h12b == _io_insn_T[9:0] ? 32'h13 : _GEN_299; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_301 = 10'h12c == _io_insn_T[9:0] ? 32'h13 : _GEN_300; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_302 = 10'h12d == _io_insn_T[9:0] ? 32'h13 : _GEN_301; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_303 = 10'h12e == _io_insn_T[9:0] ? 32'h13 : _GEN_302; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_304 = 10'h12f == _io_insn_T[9:0] ? 32'h13 : _GEN_303; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_305 = 10'h130 == _io_insn_T[9:0] ? 32'h13 : _GEN_304; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_306 = 10'h131 == _io_insn_T[9:0] ? 32'h13 : _GEN_305; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_307 = 10'h132 == _io_insn_T[9:0] ? 32'h13 : _GEN_306; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_308 = 10'h133 == _io_insn_T[9:0] ? 32'h13 : _GEN_307; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_309 = 10'h134 == _io_insn_T[9:0] ? 32'h13 : _GEN_308; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_310 = 10'h135 == _io_insn_T[9:0] ? 32'h13 : _GEN_309; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_311 = 10'h136 == _io_insn_T[9:0] ? 32'h13 : _GEN_310; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_312 = 10'h137 == _io_insn_T[9:0] ? 32'h13 : _GEN_311; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_313 = 10'h138 == _io_insn_T[9:0] ? 32'h13 : _GEN_312; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_314 = 10'h139 == _io_insn_T[9:0] ? 32'h13 : _GEN_313; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_315 = 10'h13a == _io_insn_T[9:0] ? 32'h13 : _GEN_314; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_316 = 10'h13b == _io_insn_T[9:0] ? 32'h13 : _GEN_315; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_317 = 10'h13c == _io_insn_T[9:0] ? 32'h13 : _GEN_316; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_318 = 10'h13d == _io_insn_T[9:0] ? 32'h13 : _GEN_317; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_319 = 10'h13e == _io_insn_T[9:0] ? 32'h13 : _GEN_318; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_320 = 10'h13f == _io_insn_T[9:0] ? 32'h13 : _GEN_319; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_321 = 10'h140 == _io_insn_T[9:0] ? 32'h13 : _GEN_320; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_322 = 10'h141 == _io_insn_T[9:0] ? 32'h13 : _GEN_321; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_323 = 10'h142 == _io_insn_T[9:0] ? 32'h13 : _GEN_322; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_324 = 10'h143 == _io_insn_T[9:0] ? 32'h13 : _GEN_323; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_325 = 10'h144 == _io_insn_T[9:0] ? 32'h13 : _GEN_324; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_326 = 10'h145 == _io_insn_T[9:0] ? 32'h13 : _GEN_325; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_327 = 10'h146 == _io_insn_T[9:0] ? 32'h13 : _GEN_326; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_328 = 10'h147 == _io_insn_T[9:0] ? 32'h13 : _GEN_327; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_329 = 10'h148 == _io_insn_T[9:0] ? 32'h13 : _GEN_328; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_330 = 10'h149 == _io_insn_T[9:0] ? 32'h13 : _GEN_329; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_331 = 10'h14a == _io_insn_T[9:0] ? 32'h13 : _GEN_330; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_332 = 10'h14b == _io_insn_T[9:0] ? 32'h13 : _GEN_331; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_333 = 10'h14c == _io_insn_T[9:0] ? 32'h13 : _GEN_332; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_334 = 10'h14d == _io_insn_T[9:0] ? 32'h13 : _GEN_333; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_335 = 10'h14e == _io_insn_T[9:0] ? 32'h13 : _GEN_334; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_336 = 10'h14f == _io_insn_T[9:0] ? 32'h13 : _GEN_335; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_337 = 10'h150 == _io_insn_T[9:0] ? 32'h13 : _GEN_336; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_338 = 10'h151 == _io_insn_T[9:0] ? 32'h13 : _GEN_337; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_339 = 10'h152 == _io_insn_T[9:0] ? 32'h13 : _GEN_338; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_340 = 10'h153 == _io_insn_T[9:0] ? 32'h13 : _GEN_339; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_341 = 10'h154 == _io_insn_T[9:0] ? 32'h13 : _GEN_340; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_342 = 10'h155 == _io_insn_T[9:0] ? 32'h13 : _GEN_341; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_343 = 10'h156 == _io_insn_T[9:0] ? 32'h13 : _GEN_342; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_344 = 10'h157 == _io_insn_T[9:0] ? 32'h13 : _GEN_343; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_345 = 10'h158 == _io_insn_T[9:0] ? 32'h13 : _GEN_344; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_346 = 10'h159 == _io_insn_T[9:0] ? 32'h13 : _GEN_345; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_347 = 10'h15a == _io_insn_T[9:0] ? 32'h13 : _GEN_346; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_348 = 10'h15b == _io_insn_T[9:0] ? 32'h13 : _GEN_347; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_349 = 10'h15c == _io_insn_T[9:0] ? 32'h13 : _GEN_348; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_350 = 10'h15d == _io_insn_T[9:0] ? 32'h13 : _GEN_349; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_351 = 10'h15e == _io_insn_T[9:0] ? 32'h13 : _GEN_350; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_352 = 10'h15f == _io_insn_T[9:0] ? 32'h13 : _GEN_351; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_353 = 10'h160 == _io_insn_T[9:0] ? 32'h13 : _GEN_352; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_354 = 10'h161 == _io_insn_T[9:0] ? 32'h13 : _GEN_353; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_355 = 10'h162 == _io_insn_T[9:0] ? 32'h13 : _GEN_354; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_356 = 10'h163 == _io_insn_T[9:0] ? 32'h13 : _GEN_355; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_357 = 10'h164 == _io_insn_T[9:0] ? 32'h13 : _GEN_356; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_358 = 10'h165 == _io_insn_T[9:0] ? 32'h13 : _GEN_357; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_359 = 10'h166 == _io_insn_T[9:0] ? 32'h13 : _GEN_358; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_360 = 10'h167 == _io_insn_T[9:0] ? 32'h13 : _GEN_359; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_361 = 10'h168 == _io_insn_T[9:0] ? 32'h13 : _GEN_360; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_362 = 10'h169 == _io_insn_T[9:0] ? 32'h13 : _GEN_361; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_363 = 10'h16a == _io_insn_T[9:0] ? 32'h13 : _GEN_362; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_364 = 10'h16b == _io_insn_T[9:0] ? 32'h13 : _GEN_363; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_365 = 10'h16c == _io_insn_T[9:0] ? 32'h13 : _GEN_364; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_366 = 10'h16d == _io_insn_T[9:0] ? 32'h13 : _GEN_365; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_367 = 10'h16e == _io_insn_T[9:0] ? 32'h13 : _GEN_366; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_368 = 10'h16f == _io_insn_T[9:0] ? 32'h13 : _GEN_367; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_369 = 10'h170 == _io_insn_T[9:0] ? 32'h13 : _GEN_368; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_370 = 10'h171 == _io_insn_T[9:0] ? 32'h13 : _GEN_369; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_371 = 10'h172 == _io_insn_T[9:0] ? 32'h13 : _GEN_370; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_372 = 10'h173 == _io_insn_T[9:0] ? 32'h13 : _GEN_371; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_373 = 10'h174 == _io_insn_T[9:0] ? 32'h13 : _GEN_372; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_374 = 10'h175 == _io_insn_T[9:0] ? 32'h13 : _GEN_373; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_375 = 10'h176 == _io_insn_T[9:0] ? 32'h13 : _GEN_374; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_376 = 10'h177 == _io_insn_T[9:0] ? 32'h13 : _GEN_375; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_377 = 10'h178 == _io_insn_T[9:0] ? 32'h13 : _GEN_376; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_378 = 10'h179 == _io_insn_T[9:0] ? 32'h13 : _GEN_377; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_379 = 10'h17a == _io_insn_T[9:0] ? 32'h13 : _GEN_378; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_380 = 10'h17b == _io_insn_T[9:0] ? 32'h13 : _GEN_379; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_381 = 10'h17c == _io_insn_T[9:0] ? 32'h13 : _GEN_380; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_382 = 10'h17d == _io_insn_T[9:0] ? 32'h13 : _GEN_381; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_383 = 10'h17e == _io_insn_T[9:0] ? 32'h13 : _GEN_382; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_384 = 10'h17f == _io_insn_T[9:0] ? 32'h13 : _GEN_383; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_385 = 10'h180 == _io_insn_T[9:0] ? 32'h13 : _GEN_384; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_386 = 10'h181 == _io_insn_T[9:0] ? 32'h13 : _GEN_385; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_387 = 10'h182 == _io_insn_T[9:0] ? 32'h13 : _GEN_386; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_388 = 10'h183 == _io_insn_T[9:0] ? 32'h13 : _GEN_387; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_389 = 10'h184 == _io_insn_T[9:0] ? 32'h13 : _GEN_388; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_390 = 10'h185 == _io_insn_T[9:0] ? 32'h13 : _GEN_389; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_391 = 10'h186 == _io_insn_T[9:0] ? 32'h13 : _GEN_390; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_392 = 10'h187 == _io_insn_T[9:0] ? 32'h13 : _GEN_391; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_393 = 10'h188 == _io_insn_T[9:0] ? 32'h13 : _GEN_392; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_394 = 10'h189 == _io_insn_T[9:0] ? 32'h13 : _GEN_393; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_395 = 10'h18a == _io_insn_T[9:0] ? 32'h13 : _GEN_394; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_396 = 10'h18b == _io_insn_T[9:0] ? 32'h13 : _GEN_395; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_397 = 10'h18c == _io_insn_T[9:0] ? 32'h13 : _GEN_396; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_398 = 10'h18d == _io_insn_T[9:0] ? 32'h13 : _GEN_397; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_399 = 10'h18e == _io_insn_T[9:0] ? 32'h13 : _GEN_398; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_400 = 10'h18f == _io_insn_T[9:0] ? 32'h13 : _GEN_399; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_401 = 10'h190 == _io_insn_T[9:0] ? 32'h13 : _GEN_400; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_402 = 10'h191 == _io_insn_T[9:0] ? 32'h13 : _GEN_401; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_403 = 10'h192 == _io_insn_T[9:0] ? 32'h13 : _GEN_402; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_404 = 10'h193 == _io_insn_T[9:0] ? 32'h13 : _GEN_403; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_405 = 10'h194 == _io_insn_T[9:0] ? 32'h13 : _GEN_404; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_406 = 10'h195 == _io_insn_T[9:0] ? 32'h13 : _GEN_405; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_407 = 10'h196 == _io_insn_T[9:0] ? 32'h13 : _GEN_406; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_408 = 10'h197 == _io_insn_T[9:0] ? 32'h13 : _GEN_407; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_409 = 10'h198 == _io_insn_T[9:0] ? 32'h13 : _GEN_408; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_410 = 10'h199 == _io_insn_T[9:0] ? 32'h13 : _GEN_409; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_411 = 10'h19a == _io_insn_T[9:0] ? 32'h13 : _GEN_410; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_412 = 10'h19b == _io_insn_T[9:0] ? 32'h13 : _GEN_411; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_413 = 10'h19c == _io_insn_T[9:0] ? 32'h13 : _GEN_412; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_414 = 10'h19d == _io_insn_T[9:0] ? 32'h13 : _GEN_413; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_415 = 10'h19e == _io_insn_T[9:0] ? 32'h13 : _GEN_414; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_416 = 10'h19f == _io_insn_T[9:0] ? 32'h13 : _GEN_415; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_417 = 10'h1a0 == _io_insn_T[9:0] ? 32'h13 : _GEN_416; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_418 = 10'h1a1 == _io_insn_T[9:0] ? 32'h13 : _GEN_417; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_419 = 10'h1a2 == _io_insn_T[9:0] ? 32'h13 : _GEN_418; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_420 = 10'h1a3 == _io_insn_T[9:0] ? 32'h13 : _GEN_419; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_421 = 10'h1a4 == _io_insn_T[9:0] ? 32'h13 : _GEN_420; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_422 = 10'h1a5 == _io_insn_T[9:0] ? 32'h13 : _GEN_421; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_423 = 10'h1a6 == _io_insn_T[9:0] ? 32'h13 : _GEN_422; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_424 = 10'h1a7 == _io_insn_T[9:0] ? 32'h13 : _GEN_423; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_425 = 10'h1a8 == _io_insn_T[9:0] ? 32'h13 : _GEN_424; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_426 = 10'h1a9 == _io_insn_T[9:0] ? 32'h13 : _GEN_425; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_427 = 10'h1aa == _io_insn_T[9:0] ? 32'h13 : _GEN_426; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_428 = 10'h1ab == _io_insn_T[9:0] ? 32'h13 : _GEN_427; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_429 = 10'h1ac == _io_insn_T[9:0] ? 32'h13 : _GEN_428; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_430 = 10'h1ad == _io_insn_T[9:0] ? 32'h13 : _GEN_429; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_431 = 10'h1ae == _io_insn_T[9:0] ? 32'h13 : _GEN_430; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_432 = 10'h1af == _io_insn_T[9:0] ? 32'h13 : _GEN_431; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_433 = 10'h1b0 == _io_insn_T[9:0] ? 32'h13 : _GEN_432; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_434 = 10'h1b1 == _io_insn_T[9:0] ? 32'h13 : _GEN_433; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_435 = 10'h1b2 == _io_insn_T[9:0] ? 32'h13 : _GEN_434; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_436 = 10'h1b3 == _io_insn_T[9:0] ? 32'h13 : _GEN_435; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_437 = 10'h1b4 == _io_insn_T[9:0] ? 32'h13 : _GEN_436; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_438 = 10'h1b5 == _io_insn_T[9:0] ? 32'h13 : _GEN_437; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_439 = 10'h1b6 == _io_insn_T[9:0] ? 32'h13 : _GEN_438; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_440 = 10'h1b7 == _io_insn_T[9:0] ? 32'h13 : _GEN_439; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_441 = 10'h1b8 == _io_insn_T[9:0] ? 32'h13 : _GEN_440; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_442 = 10'h1b9 == _io_insn_T[9:0] ? 32'h13 : _GEN_441; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_443 = 10'h1ba == _io_insn_T[9:0] ? 32'h13 : _GEN_442; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_444 = 10'h1bb == _io_insn_T[9:0] ? 32'h13 : _GEN_443; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_445 = 10'h1bc == _io_insn_T[9:0] ? 32'h13 : _GEN_444; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_446 = 10'h1bd == _io_insn_T[9:0] ? 32'h13 : _GEN_445; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_447 = 10'h1be == _io_insn_T[9:0] ? 32'h13 : _GEN_446; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_448 = 10'h1bf == _io_insn_T[9:0] ? 32'h13 : _GEN_447; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_449 = 10'h1c0 == _io_insn_T[9:0] ? 32'h13 : _GEN_448; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_450 = 10'h1c1 == _io_insn_T[9:0] ? 32'h13 : _GEN_449; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_451 = 10'h1c2 == _io_insn_T[9:0] ? 32'h13 : _GEN_450; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_452 = 10'h1c3 == _io_insn_T[9:0] ? 32'h13 : _GEN_451; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_453 = 10'h1c4 == _io_insn_T[9:0] ? 32'h13 : _GEN_452; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_454 = 10'h1c5 == _io_insn_T[9:0] ? 32'h13 : _GEN_453; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_455 = 10'h1c6 == _io_insn_T[9:0] ? 32'h13 : _GEN_454; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_456 = 10'h1c7 == _io_insn_T[9:0] ? 32'h13 : _GEN_455; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_457 = 10'h1c8 == _io_insn_T[9:0] ? 32'h13 : _GEN_456; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_458 = 10'h1c9 == _io_insn_T[9:0] ? 32'h13 : _GEN_457; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_459 = 10'h1ca == _io_insn_T[9:0] ? 32'h13 : _GEN_458; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_460 = 10'h1cb == _io_insn_T[9:0] ? 32'h13 : _GEN_459; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_461 = 10'h1cc == _io_insn_T[9:0] ? 32'h13 : _GEN_460; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_462 = 10'h1cd == _io_insn_T[9:0] ? 32'h13 : _GEN_461; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_463 = 10'h1ce == _io_insn_T[9:0] ? 32'h13 : _GEN_462; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_464 = 10'h1cf == _io_insn_T[9:0] ? 32'h13 : _GEN_463; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_465 = 10'h1d0 == _io_insn_T[9:0] ? 32'h13 : _GEN_464; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_466 = 10'h1d1 == _io_insn_T[9:0] ? 32'h13 : _GEN_465; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_467 = 10'h1d2 == _io_insn_T[9:0] ? 32'h13 : _GEN_466; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_468 = 10'h1d3 == _io_insn_T[9:0] ? 32'h13 : _GEN_467; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_469 = 10'h1d4 == _io_insn_T[9:0] ? 32'h13 : _GEN_468; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_470 = 10'h1d5 == _io_insn_T[9:0] ? 32'h13 : _GEN_469; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_471 = 10'h1d6 == _io_insn_T[9:0] ? 32'h13 : _GEN_470; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_472 = 10'h1d7 == _io_insn_T[9:0] ? 32'h13 : _GEN_471; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_473 = 10'h1d8 == _io_insn_T[9:0] ? 32'h13 : _GEN_472; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_474 = 10'h1d9 == _io_insn_T[9:0] ? 32'h13 : _GEN_473; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_475 = 10'h1da == _io_insn_T[9:0] ? 32'h13 : _GEN_474; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_476 = 10'h1db == _io_insn_T[9:0] ? 32'h13 : _GEN_475; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_477 = 10'h1dc == _io_insn_T[9:0] ? 32'h13 : _GEN_476; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_478 = 10'h1dd == _io_insn_T[9:0] ? 32'h13 : _GEN_477; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_479 = 10'h1de == _io_insn_T[9:0] ? 32'h13 : _GEN_478; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_480 = 10'h1df == _io_insn_T[9:0] ? 32'h13 : _GEN_479; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_481 = 10'h1e0 == _io_insn_T[9:0] ? 32'h13 : _GEN_480; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_482 = 10'h1e1 == _io_insn_T[9:0] ? 32'h13 : _GEN_481; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_483 = 10'h1e2 == _io_insn_T[9:0] ? 32'h13 : _GEN_482; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_484 = 10'h1e3 == _io_insn_T[9:0] ? 32'h13 : _GEN_483; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_485 = 10'h1e4 == _io_insn_T[9:0] ? 32'h13 : _GEN_484; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_486 = 10'h1e5 == _io_insn_T[9:0] ? 32'h13 : _GEN_485; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_487 = 10'h1e6 == _io_insn_T[9:0] ? 32'h13 : _GEN_486; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_488 = 10'h1e7 == _io_insn_T[9:0] ? 32'h13 : _GEN_487; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_489 = 10'h1e8 == _io_insn_T[9:0] ? 32'h13 : _GEN_488; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_490 = 10'h1e9 == _io_insn_T[9:0] ? 32'h13 : _GEN_489; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_491 = 10'h1ea == _io_insn_T[9:0] ? 32'h13 : _GEN_490; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_492 = 10'h1eb == _io_insn_T[9:0] ? 32'h13 : _GEN_491; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_493 = 10'h1ec == _io_insn_T[9:0] ? 32'h13 : _GEN_492; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_494 = 10'h1ed == _io_insn_T[9:0] ? 32'h13 : _GEN_493; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_495 = 10'h1ee == _io_insn_T[9:0] ? 32'h13 : _GEN_494; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_496 = 10'h1ef == _io_insn_T[9:0] ? 32'h13 : _GEN_495; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_497 = 10'h1f0 == _io_insn_T[9:0] ? 32'h13 : _GEN_496; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_498 = 10'h1f1 == _io_insn_T[9:0] ? 32'h13 : _GEN_497; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_499 = 10'h1f2 == _io_insn_T[9:0] ? 32'h13 : _GEN_498; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_500 = 10'h1f3 == _io_insn_T[9:0] ? 32'h13 : _GEN_499; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_501 = 10'h1f4 == _io_insn_T[9:0] ? 32'h13 : _GEN_500; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_502 = 10'h1f5 == _io_insn_T[9:0] ? 32'h13 : _GEN_501; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_503 = 10'h1f6 == _io_insn_T[9:0] ? 32'h13 : _GEN_502; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_504 = 10'h1f7 == _io_insn_T[9:0] ? 32'h13 : _GEN_503; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_505 = 10'h1f8 == _io_insn_T[9:0] ? 32'h13 : _GEN_504; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_506 = 10'h1f9 == _io_insn_T[9:0] ? 32'h13 : _GEN_505; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_507 = 10'h1fa == _io_insn_T[9:0] ? 32'h13 : _GEN_506; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_508 = 10'h1fb == _io_insn_T[9:0] ? 32'h13 : _GEN_507; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_509 = 10'h1fc == _io_insn_T[9:0] ? 32'h13 : _GEN_508; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_510 = 10'h1fd == _io_insn_T[9:0] ? 32'h13 : _GEN_509; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_511 = 10'h1fe == _io_insn_T[9:0] ? 32'h13 : _GEN_510; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_512 = 10'h1ff == _io_insn_T[9:0] ? 32'h13 : _GEN_511; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_513 = 10'h200 == _io_insn_T[9:0] ? 32'h13 : _GEN_512; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_514 = 10'h201 == _io_insn_T[9:0] ? 32'h13 : _GEN_513; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_515 = 10'h202 == _io_insn_T[9:0] ? 32'h13 : _GEN_514; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_516 = 10'h203 == _io_insn_T[9:0] ? 32'h13 : _GEN_515; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_517 = 10'h204 == _io_insn_T[9:0] ? 32'h13 : _GEN_516; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_518 = 10'h205 == _io_insn_T[9:0] ? 32'h13 : _GEN_517; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_519 = 10'h206 == _io_insn_T[9:0] ? 32'h13 : _GEN_518; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_520 = 10'h207 == _io_insn_T[9:0] ? 32'h13 : _GEN_519; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_521 = 10'h208 == _io_insn_T[9:0] ? 32'h13 : _GEN_520; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_522 = 10'h209 == _io_insn_T[9:0] ? 32'h13 : _GEN_521; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_523 = 10'h20a == _io_insn_T[9:0] ? 32'h13 : _GEN_522; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_524 = 10'h20b == _io_insn_T[9:0] ? 32'h13 : _GEN_523; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_525 = 10'h20c == _io_insn_T[9:0] ? 32'h13 : _GEN_524; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_526 = 10'h20d == _io_insn_T[9:0] ? 32'h13 : _GEN_525; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_527 = 10'h20e == _io_insn_T[9:0] ? 32'h13 : _GEN_526; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_528 = 10'h20f == _io_insn_T[9:0] ? 32'h13 : _GEN_527; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_529 = 10'h210 == _io_insn_T[9:0] ? 32'h13 : _GEN_528; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_530 = 10'h211 == _io_insn_T[9:0] ? 32'h13 : _GEN_529; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_531 = 10'h212 == _io_insn_T[9:0] ? 32'h13 : _GEN_530; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_532 = 10'h213 == _io_insn_T[9:0] ? 32'h13 : _GEN_531; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_533 = 10'h214 == _io_insn_T[9:0] ? 32'h13 : _GEN_532; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_534 = 10'h215 == _io_insn_T[9:0] ? 32'h13 : _GEN_533; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_535 = 10'h216 == _io_insn_T[9:0] ? 32'h13 : _GEN_534; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_536 = 10'h217 == _io_insn_T[9:0] ? 32'h13 : _GEN_535; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_537 = 10'h218 == _io_insn_T[9:0] ? 32'h13 : _GEN_536; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_538 = 10'h219 == _io_insn_T[9:0] ? 32'h13 : _GEN_537; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_539 = 10'h21a == _io_insn_T[9:0] ? 32'h13 : _GEN_538; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_540 = 10'h21b == _io_insn_T[9:0] ? 32'h13 : _GEN_539; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_541 = 10'h21c == _io_insn_T[9:0] ? 32'h13 : _GEN_540; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_542 = 10'h21d == _io_insn_T[9:0] ? 32'h13 : _GEN_541; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_543 = 10'h21e == _io_insn_T[9:0] ? 32'h13 : _GEN_542; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_544 = 10'h21f == _io_insn_T[9:0] ? 32'h13 : _GEN_543; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_545 = 10'h220 == _io_insn_T[9:0] ? 32'h13 : _GEN_544; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_546 = 10'h221 == _io_insn_T[9:0] ? 32'h13 : _GEN_545; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_547 = 10'h222 == _io_insn_T[9:0] ? 32'h13 : _GEN_546; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_548 = 10'h223 == _io_insn_T[9:0] ? 32'h13 : _GEN_547; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_549 = 10'h224 == _io_insn_T[9:0] ? 32'h13 : _GEN_548; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_550 = 10'h225 == _io_insn_T[9:0] ? 32'h13 : _GEN_549; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_551 = 10'h226 == _io_insn_T[9:0] ? 32'h13 : _GEN_550; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_552 = 10'h227 == _io_insn_T[9:0] ? 32'h13 : _GEN_551; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_553 = 10'h228 == _io_insn_T[9:0] ? 32'h13 : _GEN_552; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_554 = 10'h229 == _io_insn_T[9:0] ? 32'h13 : _GEN_553; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_555 = 10'h22a == _io_insn_T[9:0] ? 32'h13 : _GEN_554; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_556 = 10'h22b == _io_insn_T[9:0] ? 32'h13 : _GEN_555; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_557 = 10'h22c == _io_insn_T[9:0] ? 32'h13 : _GEN_556; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_558 = 10'h22d == _io_insn_T[9:0] ? 32'h13 : _GEN_557; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_559 = 10'h22e == _io_insn_T[9:0] ? 32'h13 : _GEN_558; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_560 = 10'h22f == _io_insn_T[9:0] ? 32'h13 : _GEN_559; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_561 = 10'h230 == _io_insn_T[9:0] ? 32'h13 : _GEN_560; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_562 = 10'h231 == _io_insn_T[9:0] ? 32'h13 : _GEN_561; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_563 = 10'h232 == _io_insn_T[9:0] ? 32'h13 : _GEN_562; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_564 = 10'h233 == _io_insn_T[9:0] ? 32'h13 : _GEN_563; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_565 = 10'h234 == _io_insn_T[9:0] ? 32'h13 : _GEN_564; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_566 = 10'h235 == _io_insn_T[9:0] ? 32'h13 : _GEN_565; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_567 = 10'h236 == _io_insn_T[9:0] ? 32'h13 : _GEN_566; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_568 = 10'h237 == _io_insn_T[9:0] ? 32'h13 : _GEN_567; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_569 = 10'h238 == _io_insn_T[9:0] ? 32'h13 : _GEN_568; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_570 = 10'h239 == _io_insn_T[9:0] ? 32'h13 : _GEN_569; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_571 = 10'h23a == _io_insn_T[9:0] ? 32'h13 : _GEN_570; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_572 = 10'h23b == _io_insn_T[9:0] ? 32'h13 : _GEN_571; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_573 = 10'h23c == _io_insn_T[9:0] ? 32'h13 : _GEN_572; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_574 = 10'h23d == _io_insn_T[9:0] ? 32'h13 : _GEN_573; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_575 = 10'h23e == _io_insn_T[9:0] ? 32'h13 : _GEN_574; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_576 = 10'h23f == _io_insn_T[9:0] ? 32'h13 : _GEN_575; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_577 = 10'h240 == _io_insn_T[9:0] ? 32'h13 : _GEN_576; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_578 = 10'h241 == _io_insn_T[9:0] ? 32'h13 : _GEN_577; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_579 = 10'h242 == _io_insn_T[9:0] ? 32'h13 : _GEN_578; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_580 = 10'h243 == _io_insn_T[9:0] ? 32'h13 : _GEN_579; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_581 = 10'h244 == _io_insn_T[9:0] ? 32'h13 : _GEN_580; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_582 = 10'h245 == _io_insn_T[9:0] ? 32'h13 : _GEN_581; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_583 = 10'h246 == _io_insn_T[9:0] ? 32'h13 : _GEN_582; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_584 = 10'h247 == _io_insn_T[9:0] ? 32'h13 : _GEN_583; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_585 = 10'h248 == _io_insn_T[9:0] ? 32'h13 : _GEN_584; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_586 = 10'h249 == _io_insn_T[9:0] ? 32'h13 : _GEN_585; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_587 = 10'h24a == _io_insn_T[9:0] ? 32'h13 : _GEN_586; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_588 = 10'h24b == _io_insn_T[9:0] ? 32'h13 : _GEN_587; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_589 = 10'h24c == _io_insn_T[9:0] ? 32'h13 : _GEN_588; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_590 = 10'h24d == _io_insn_T[9:0] ? 32'h13 : _GEN_589; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_591 = 10'h24e == _io_insn_T[9:0] ? 32'h13 : _GEN_590; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_592 = 10'h24f == _io_insn_T[9:0] ? 32'h13 : _GEN_591; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_593 = 10'h250 == _io_insn_T[9:0] ? 32'h13 : _GEN_592; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_594 = 10'h251 == _io_insn_T[9:0] ? 32'h13 : _GEN_593; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_595 = 10'h252 == _io_insn_T[9:0] ? 32'h13 : _GEN_594; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_596 = 10'h253 == _io_insn_T[9:0] ? 32'h13 : _GEN_595; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_597 = 10'h254 == _io_insn_T[9:0] ? 32'h13 : _GEN_596; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_598 = 10'h255 == _io_insn_T[9:0] ? 32'h13 : _GEN_597; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_599 = 10'h256 == _io_insn_T[9:0] ? 32'h13 : _GEN_598; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_600 = 10'h257 == _io_insn_T[9:0] ? 32'h13 : _GEN_599; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_601 = 10'h258 == _io_insn_T[9:0] ? 32'h13 : _GEN_600; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_602 = 10'h259 == _io_insn_T[9:0] ? 32'h13 : _GEN_601; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_603 = 10'h25a == _io_insn_T[9:0] ? 32'h13 : _GEN_602; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_604 = 10'h25b == _io_insn_T[9:0] ? 32'h13 : _GEN_603; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_605 = 10'h25c == _io_insn_T[9:0] ? 32'h13 : _GEN_604; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_606 = 10'h25d == _io_insn_T[9:0] ? 32'h13 : _GEN_605; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_607 = 10'h25e == _io_insn_T[9:0] ? 32'h13 : _GEN_606; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_608 = 10'h25f == _io_insn_T[9:0] ? 32'h13 : _GEN_607; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_609 = 10'h260 == _io_insn_T[9:0] ? 32'h13 : _GEN_608; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_610 = 10'h261 == _io_insn_T[9:0] ? 32'h13 : _GEN_609; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_611 = 10'h262 == _io_insn_T[9:0] ? 32'h13 : _GEN_610; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_612 = 10'h263 == _io_insn_T[9:0] ? 32'h13 : _GEN_611; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_613 = 10'h264 == _io_insn_T[9:0] ? 32'h13 : _GEN_612; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_614 = 10'h265 == _io_insn_T[9:0] ? 32'h13 : _GEN_613; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_615 = 10'h266 == _io_insn_T[9:0] ? 32'h13 : _GEN_614; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_616 = 10'h267 == _io_insn_T[9:0] ? 32'h13 : _GEN_615; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_617 = 10'h268 == _io_insn_T[9:0] ? 32'h13 : _GEN_616; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_618 = 10'h269 == _io_insn_T[9:0] ? 32'h13 : _GEN_617; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_619 = 10'h26a == _io_insn_T[9:0] ? 32'h13 : _GEN_618; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_620 = 10'h26b == _io_insn_T[9:0] ? 32'h13 : _GEN_619; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_621 = 10'h26c == _io_insn_T[9:0] ? 32'h13 : _GEN_620; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_622 = 10'h26d == _io_insn_T[9:0] ? 32'h13 : _GEN_621; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_623 = 10'h26e == _io_insn_T[9:0] ? 32'h13 : _GEN_622; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_624 = 10'h26f == _io_insn_T[9:0] ? 32'h13 : _GEN_623; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_625 = 10'h270 == _io_insn_T[9:0] ? 32'h13 : _GEN_624; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_626 = 10'h271 == _io_insn_T[9:0] ? 32'h13 : _GEN_625; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_627 = 10'h272 == _io_insn_T[9:0] ? 32'h13 : _GEN_626; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_628 = 10'h273 == _io_insn_T[9:0] ? 32'h13 : _GEN_627; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_629 = 10'h274 == _io_insn_T[9:0] ? 32'h13 : _GEN_628; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_630 = 10'h275 == _io_insn_T[9:0] ? 32'h13 : _GEN_629; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_631 = 10'h276 == _io_insn_T[9:0] ? 32'h13 : _GEN_630; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_632 = 10'h277 == _io_insn_T[9:0] ? 32'h13 : _GEN_631; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_633 = 10'h278 == _io_insn_T[9:0] ? 32'h13 : _GEN_632; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_634 = 10'h279 == _io_insn_T[9:0] ? 32'h13 : _GEN_633; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_635 = 10'h27a == _io_insn_T[9:0] ? 32'h13 : _GEN_634; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_636 = 10'h27b == _io_insn_T[9:0] ? 32'h13 : _GEN_635; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_637 = 10'h27c == _io_insn_T[9:0] ? 32'h13 : _GEN_636; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_638 = 10'h27d == _io_insn_T[9:0] ? 32'h13 : _GEN_637; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_639 = 10'h27e == _io_insn_T[9:0] ? 32'h13 : _GEN_638; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_640 = 10'h27f == _io_insn_T[9:0] ? 32'h13 : _GEN_639; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_641 = 10'h280 == _io_insn_T[9:0] ? 32'h13 : _GEN_640; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_642 = 10'h281 == _io_insn_T[9:0] ? 32'h13 : _GEN_641; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_643 = 10'h282 == _io_insn_T[9:0] ? 32'h13 : _GEN_642; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_644 = 10'h283 == _io_insn_T[9:0] ? 32'h13 : _GEN_643; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_645 = 10'h284 == _io_insn_T[9:0] ? 32'h13 : _GEN_644; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_646 = 10'h285 == _io_insn_T[9:0] ? 32'h13 : _GEN_645; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_647 = 10'h286 == _io_insn_T[9:0] ? 32'h13 : _GEN_646; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_648 = 10'h287 == _io_insn_T[9:0] ? 32'h13 : _GEN_647; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_649 = 10'h288 == _io_insn_T[9:0] ? 32'h13 : _GEN_648; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_650 = 10'h289 == _io_insn_T[9:0] ? 32'h13 : _GEN_649; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_651 = 10'h28a == _io_insn_T[9:0] ? 32'h13 : _GEN_650; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_652 = 10'h28b == _io_insn_T[9:0] ? 32'h13 : _GEN_651; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_653 = 10'h28c == _io_insn_T[9:0] ? 32'h13 : _GEN_652; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_654 = 10'h28d == _io_insn_T[9:0] ? 32'h13 : _GEN_653; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_655 = 10'h28e == _io_insn_T[9:0] ? 32'h13 : _GEN_654; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_656 = 10'h28f == _io_insn_T[9:0] ? 32'h13 : _GEN_655; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_657 = 10'h290 == _io_insn_T[9:0] ? 32'h13 : _GEN_656; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_658 = 10'h291 == _io_insn_T[9:0] ? 32'h13 : _GEN_657; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_659 = 10'h292 == _io_insn_T[9:0] ? 32'h13 : _GEN_658; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_660 = 10'h293 == _io_insn_T[9:0] ? 32'h13 : _GEN_659; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_661 = 10'h294 == _io_insn_T[9:0] ? 32'h13 : _GEN_660; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_662 = 10'h295 == _io_insn_T[9:0] ? 32'h13 : _GEN_661; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_663 = 10'h296 == _io_insn_T[9:0] ? 32'h13 : _GEN_662; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_664 = 10'h297 == _io_insn_T[9:0] ? 32'h13 : _GEN_663; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_665 = 10'h298 == _io_insn_T[9:0] ? 32'h13 : _GEN_664; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_666 = 10'h299 == _io_insn_T[9:0] ? 32'h13 : _GEN_665; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_667 = 10'h29a == _io_insn_T[9:0] ? 32'h13 : _GEN_666; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_668 = 10'h29b == _io_insn_T[9:0] ? 32'h13 : _GEN_667; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_669 = 10'h29c == _io_insn_T[9:0] ? 32'h13 : _GEN_668; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_670 = 10'h29d == _io_insn_T[9:0] ? 32'h13 : _GEN_669; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_671 = 10'h29e == _io_insn_T[9:0] ? 32'h13 : _GEN_670; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_672 = 10'h29f == _io_insn_T[9:0] ? 32'h13 : _GEN_671; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_673 = 10'h2a0 == _io_insn_T[9:0] ? 32'h13 : _GEN_672; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_674 = 10'h2a1 == _io_insn_T[9:0] ? 32'h13 : _GEN_673; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_675 = 10'h2a2 == _io_insn_T[9:0] ? 32'h13 : _GEN_674; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_676 = 10'h2a3 == _io_insn_T[9:0] ? 32'h13 : _GEN_675; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_677 = 10'h2a4 == _io_insn_T[9:0] ? 32'h13 : _GEN_676; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_678 = 10'h2a5 == _io_insn_T[9:0] ? 32'h13 : _GEN_677; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_679 = 10'h2a6 == _io_insn_T[9:0] ? 32'h13 : _GEN_678; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_680 = 10'h2a7 == _io_insn_T[9:0] ? 32'h13 : _GEN_679; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_681 = 10'h2a8 == _io_insn_T[9:0] ? 32'h13 : _GEN_680; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_682 = 10'h2a9 == _io_insn_T[9:0] ? 32'h13 : _GEN_681; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_683 = 10'h2aa == _io_insn_T[9:0] ? 32'h13 : _GEN_682; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_684 = 10'h2ab == _io_insn_T[9:0] ? 32'h13 : _GEN_683; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_685 = 10'h2ac == _io_insn_T[9:0] ? 32'h13 : _GEN_684; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_686 = 10'h2ad == _io_insn_T[9:0] ? 32'h13 : _GEN_685; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_687 = 10'h2ae == _io_insn_T[9:0] ? 32'h13 : _GEN_686; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_688 = 10'h2af == _io_insn_T[9:0] ? 32'h13 : _GEN_687; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_689 = 10'h2b0 == _io_insn_T[9:0] ? 32'h13 : _GEN_688; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_690 = 10'h2b1 == _io_insn_T[9:0] ? 32'h13 : _GEN_689; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_691 = 10'h2b2 == _io_insn_T[9:0] ? 32'h13 : _GEN_690; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_692 = 10'h2b3 == _io_insn_T[9:0] ? 32'h13 : _GEN_691; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_693 = 10'h2b4 == _io_insn_T[9:0] ? 32'h13 : _GEN_692; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_694 = 10'h2b5 == _io_insn_T[9:0] ? 32'h13 : _GEN_693; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_695 = 10'h2b6 == _io_insn_T[9:0] ? 32'h13 : _GEN_694; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_696 = 10'h2b7 == _io_insn_T[9:0] ? 32'h13 : _GEN_695; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_697 = 10'h2b8 == _io_insn_T[9:0] ? 32'h13 : _GEN_696; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_698 = 10'h2b9 == _io_insn_T[9:0] ? 32'h13 : _GEN_697; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_699 = 10'h2ba == _io_insn_T[9:0] ? 32'h13 : _GEN_698; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_700 = 10'h2bb == _io_insn_T[9:0] ? 32'h13 : _GEN_699; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_701 = 10'h2bc == _io_insn_T[9:0] ? 32'h13 : _GEN_700; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_702 = 10'h2bd == _io_insn_T[9:0] ? 32'h13 : _GEN_701; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_703 = 10'h2be == _io_insn_T[9:0] ? 32'h13 : _GEN_702; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_704 = 10'h2bf == _io_insn_T[9:0] ? 32'h13 : _GEN_703; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_705 = 10'h2c0 == _io_insn_T[9:0] ? 32'h13 : _GEN_704; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_706 = 10'h2c1 == _io_insn_T[9:0] ? 32'h13 : _GEN_705; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_707 = 10'h2c2 == _io_insn_T[9:0] ? 32'h13 : _GEN_706; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_708 = 10'h2c3 == _io_insn_T[9:0] ? 32'h13 : _GEN_707; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_709 = 10'h2c4 == _io_insn_T[9:0] ? 32'h13 : _GEN_708; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_710 = 10'h2c5 == _io_insn_T[9:0] ? 32'h13 : _GEN_709; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_711 = 10'h2c6 == _io_insn_T[9:0] ? 32'h13 : _GEN_710; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_712 = 10'h2c7 == _io_insn_T[9:0] ? 32'h13 : _GEN_711; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_713 = 10'h2c8 == _io_insn_T[9:0] ? 32'h13 : _GEN_712; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_714 = 10'h2c9 == _io_insn_T[9:0] ? 32'h13 : _GEN_713; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_715 = 10'h2ca == _io_insn_T[9:0] ? 32'h13 : _GEN_714; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_716 = 10'h2cb == _io_insn_T[9:0] ? 32'h13 : _GEN_715; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_717 = 10'h2cc == _io_insn_T[9:0] ? 32'h13 : _GEN_716; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_718 = 10'h2cd == _io_insn_T[9:0] ? 32'h13 : _GEN_717; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_719 = 10'h2ce == _io_insn_T[9:0] ? 32'h13 : _GEN_718; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_720 = 10'h2cf == _io_insn_T[9:0] ? 32'h13 : _GEN_719; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_721 = 10'h2d0 == _io_insn_T[9:0] ? 32'h13 : _GEN_720; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_722 = 10'h2d1 == _io_insn_T[9:0] ? 32'h13 : _GEN_721; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_723 = 10'h2d2 == _io_insn_T[9:0] ? 32'h13 : _GEN_722; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_724 = 10'h2d3 == _io_insn_T[9:0] ? 32'h13 : _GEN_723; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_725 = 10'h2d4 == _io_insn_T[9:0] ? 32'h13 : _GEN_724; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_726 = 10'h2d5 == _io_insn_T[9:0] ? 32'h13 : _GEN_725; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_727 = 10'h2d6 == _io_insn_T[9:0] ? 32'h13 : _GEN_726; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_728 = 10'h2d7 == _io_insn_T[9:0] ? 32'h13 : _GEN_727; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_729 = 10'h2d8 == _io_insn_T[9:0] ? 32'h13 : _GEN_728; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_730 = 10'h2d9 == _io_insn_T[9:0] ? 32'h13 : _GEN_729; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_731 = 10'h2da == _io_insn_T[9:0] ? 32'h13 : _GEN_730; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_732 = 10'h2db == _io_insn_T[9:0] ? 32'h13 : _GEN_731; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_733 = 10'h2dc == _io_insn_T[9:0] ? 32'h13 : _GEN_732; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_734 = 10'h2dd == _io_insn_T[9:0] ? 32'h13 : _GEN_733; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_735 = 10'h2de == _io_insn_T[9:0] ? 32'h13 : _GEN_734; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_736 = 10'h2df == _io_insn_T[9:0] ? 32'h13 : _GEN_735; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_737 = 10'h2e0 == _io_insn_T[9:0] ? 32'h13 : _GEN_736; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_738 = 10'h2e1 == _io_insn_T[9:0] ? 32'h13 : _GEN_737; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_739 = 10'h2e2 == _io_insn_T[9:0] ? 32'h13 : _GEN_738; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_740 = 10'h2e3 == _io_insn_T[9:0] ? 32'h13 : _GEN_739; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_741 = 10'h2e4 == _io_insn_T[9:0] ? 32'h13 : _GEN_740; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_742 = 10'h2e5 == _io_insn_T[9:0] ? 32'h13 : _GEN_741; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_743 = 10'h2e6 == _io_insn_T[9:0] ? 32'h13 : _GEN_742; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_744 = 10'h2e7 == _io_insn_T[9:0] ? 32'h13 : _GEN_743; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_745 = 10'h2e8 == _io_insn_T[9:0] ? 32'h13 : _GEN_744; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_746 = 10'h2e9 == _io_insn_T[9:0] ? 32'h13 : _GEN_745; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_747 = 10'h2ea == _io_insn_T[9:0] ? 32'h13 : _GEN_746; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_748 = 10'h2eb == _io_insn_T[9:0] ? 32'h13 : _GEN_747; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_749 = 10'h2ec == _io_insn_T[9:0] ? 32'h13 : _GEN_748; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_750 = 10'h2ed == _io_insn_T[9:0] ? 32'h13 : _GEN_749; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_751 = 10'h2ee == _io_insn_T[9:0] ? 32'h13 : _GEN_750; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_752 = 10'h2ef == _io_insn_T[9:0] ? 32'h13 : _GEN_751; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_753 = 10'h2f0 == _io_insn_T[9:0] ? 32'h13 : _GEN_752; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_754 = 10'h2f1 == _io_insn_T[9:0] ? 32'h13 : _GEN_753; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_755 = 10'h2f2 == _io_insn_T[9:0] ? 32'h13 : _GEN_754; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_756 = 10'h2f3 == _io_insn_T[9:0] ? 32'h13 : _GEN_755; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_757 = 10'h2f4 == _io_insn_T[9:0] ? 32'h13 : _GEN_756; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_758 = 10'h2f5 == _io_insn_T[9:0] ? 32'h13 : _GEN_757; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_759 = 10'h2f6 == _io_insn_T[9:0] ? 32'h13 : _GEN_758; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_760 = 10'h2f7 == _io_insn_T[9:0] ? 32'h13 : _GEN_759; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_761 = 10'h2f8 == _io_insn_T[9:0] ? 32'h13 : _GEN_760; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_762 = 10'h2f9 == _io_insn_T[9:0] ? 32'h13 : _GEN_761; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_763 = 10'h2fa == _io_insn_T[9:0] ? 32'h13 : _GEN_762; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_764 = 10'h2fb == _io_insn_T[9:0] ? 32'h13 : _GEN_763; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_765 = 10'h2fc == _io_insn_T[9:0] ? 32'h13 : _GEN_764; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_766 = 10'h2fd == _io_insn_T[9:0] ? 32'h13 : _GEN_765; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_767 = 10'h2fe == _io_insn_T[9:0] ? 32'h13 : _GEN_766; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_768 = 10'h2ff == _io_insn_T[9:0] ? 32'h13 : _GEN_767; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_769 = 10'h300 == _io_insn_T[9:0] ? 32'h13 : _GEN_768; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_770 = 10'h301 == _io_insn_T[9:0] ? 32'h13 : _GEN_769; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_771 = 10'h302 == _io_insn_T[9:0] ? 32'h13 : _GEN_770; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_772 = 10'h303 == _io_insn_T[9:0] ? 32'h13 : _GEN_771; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_773 = 10'h304 == _io_insn_T[9:0] ? 32'h13 : _GEN_772; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_774 = 10'h305 == _io_insn_T[9:0] ? 32'h13 : _GEN_773; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_775 = 10'h306 == _io_insn_T[9:0] ? 32'h13 : _GEN_774; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_776 = 10'h307 == _io_insn_T[9:0] ? 32'h13 : _GEN_775; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_777 = 10'h308 == _io_insn_T[9:0] ? 32'h13 : _GEN_776; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_778 = 10'h309 == _io_insn_T[9:0] ? 32'h13 : _GEN_777; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_779 = 10'h30a == _io_insn_T[9:0] ? 32'h13 : _GEN_778; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_780 = 10'h30b == _io_insn_T[9:0] ? 32'h13 : _GEN_779; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_781 = 10'h30c == _io_insn_T[9:0] ? 32'h13 : _GEN_780; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_782 = 10'h30d == _io_insn_T[9:0] ? 32'h13 : _GEN_781; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_783 = 10'h30e == _io_insn_T[9:0] ? 32'h13 : _GEN_782; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_784 = 10'h30f == _io_insn_T[9:0] ? 32'h13 : _GEN_783; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_785 = 10'h310 == _io_insn_T[9:0] ? 32'h13 : _GEN_784; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_786 = 10'h311 == _io_insn_T[9:0] ? 32'h13 : _GEN_785; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_787 = 10'h312 == _io_insn_T[9:0] ? 32'h13 : _GEN_786; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_788 = 10'h313 == _io_insn_T[9:0] ? 32'h13 : _GEN_787; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_789 = 10'h314 == _io_insn_T[9:0] ? 32'h13 : _GEN_788; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_790 = 10'h315 == _io_insn_T[9:0] ? 32'h13 : _GEN_789; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_791 = 10'h316 == _io_insn_T[9:0] ? 32'h13 : _GEN_790; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_792 = 10'h317 == _io_insn_T[9:0] ? 32'h13 : _GEN_791; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_793 = 10'h318 == _io_insn_T[9:0] ? 32'h13 : _GEN_792; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_794 = 10'h319 == _io_insn_T[9:0] ? 32'h13 : _GEN_793; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_795 = 10'h31a == _io_insn_T[9:0] ? 32'h13 : _GEN_794; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_796 = 10'h31b == _io_insn_T[9:0] ? 32'h13 : _GEN_795; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_797 = 10'h31c == _io_insn_T[9:0] ? 32'h13 : _GEN_796; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_798 = 10'h31d == _io_insn_T[9:0] ? 32'h13 : _GEN_797; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_799 = 10'h31e == _io_insn_T[9:0] ? 32'h13 : _GEN_798; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_800 = 10'h31f == _io_insn_T[9:0] ? 32'h13 : _GEN_799; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_801 = 10'h320 == _io_insn_T[9:0] ? 32'h13 : _GEN_800; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_802 = 10'h321 == _io_insn_T[9:0] ? 32'h13 : _GEN_801; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_803 = 10'h322 == _io_insn_T[9:0] ? 32'h13 : _GEN_802; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_804 = 10'h323 == _io_insn_T[9:0] ? 32'h13 : _GEN_803; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_805 = 10'h324 == _io_insn_T[9:0] ? 32'h13 : _GEN_804; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_806 = 10'h325 == _io_insn_T[9:0] ? 32'h13 : _GEN_805; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_807 = 10'h326 == _io_insn_T[9:0] ? 32'h13 : _GEN_806; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_808 = 10'h327 == _io_insn_T[9:0] ? 32'h13 : _GEN_807; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_809 = 10'h328 == _io_insn_T[9:0] ? 32'h13 : _GEN_808; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_810 = 10'h329 == _io_insn_T[9:0] ? 32'h13 : _GEN_809; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_811 = 10'h32a == _io_insn_T[9:0] ? 32'h13 : _GEN_810; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_812 = 10'h32b == _io_insn_T[9:0] ? 32'h13 : _GEN_811; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_813 = 10'h32c == _io_insn_T[9:0] ? 32'h13 : _GEN_812; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_814 = 10'h32d == _io_insn_T[9:0] ? 32'h13 : _GEN_813; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_815 = 10'h32e == _io_insn_T[9:0] ? 32'h13 : _GEN_814; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_816 = 10'h32f == _io_insn_T[9:0] ? 32'h13 : _GEN_815; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_817 = 10'h330 == _io_insn_T[9:0] ? 32'h13 : _GEN_816; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_818 = 10'h331 == _io_insn_T[9:0] ? 32'h13 : _GEN_817; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_819 = 10'h332 == _io_insn_T[9:0] ? 32'h13 : _GEN_818; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_820 = 10'h333 == _io_insn_T[9:0] ? 32'h13 : _GEN_819; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_821 = 10'h334 == _io_insn_T[9:0] ? 32'h13 : _GEN_820; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_822 = 10'h335 == _io_insn_T[9:0] ? 32'h13 : _GEN_821; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_823 = 10'h336 == _io_insn_T[9:0] ? 32'h13 : _GEN_822; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_824 = 10'h337 == _io_insn_T[9:0] ? 32'h13 : _GEN_823; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_825 = 10'h338 == _io_insn_T[9:0] ? 32'h13 : _GEN_824; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_826 = 10'h339 == _io_insn_T[9:0] ? 32'h13 : _GEN_825; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_827 = 10'h33a == _io_insn_T[9:0] ? 32'h13 : _GEN_826; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_828 = 10'h33b == _io_insn_T[9:0] ? 32'h13 : _GEN_827; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_829 = 10'h33c == _io_insn_T[9:0] ? 32'h13 : _GEN_828; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_830 = 10'h33d == _io_insn_T[9:0] ? 32'h13 : _GEN_829; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_831 = 10'h33e == _io_insn_T[9:0] ? 32'h13 : _GEN_830; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_832 = 10'h33f == _io_insn_T[9:0] ? 32'h13 : _GEN_831; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_833 = 10'h340 == _io_insn_T[9:0] ? 32'h13 : _GEN_832; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_834 = 10'h341 == _io_insn_T[9:0] ? 32'h13 : _GEN_833; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_835 = 10'h342 == _io_insn_T[9:0] ? 32'h13 : _GEN_834; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_836 = 10'h343 == _io_insn_T[9:0] ? 32'h13 : _GEN_835; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_837 = 10'h344 == _io_insn_T[9:0] ? 32'h13 : _GEN_836; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_838 = 10'h345 == _io_insn_T[9:0] ? 32'h13 : _GEN_837; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_839 = 10'h346 == _io_insn_T[9:0] ? 32'h13 : _GEN_838; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_840 = 10'h347 == _io_insn_T[9:0] ? 32'h13 : _GEN_839; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_841 = 10'h348 == _io_insn_T[9:0] ? 32'h13 : _GEN_840; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_842 = 10'h349 == _io_insn_T[9:0] ? 32'h13 : _GEN_841; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_843 = 10'h34a == _io_insn_T[9:0] ? 32'h13 : _GEN_842; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_844 = 10'h34b == _io_insn_T[9:0] ? 32'h13 : _GEN_843; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_845 = 10'h34c == _io_insn_T[9:0] ? 32'h13 : _GEN_844; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_846 = 10'h34d == _io_insn_T[9:0] ? 32'h13 : _GEN_845; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_847 = 10'h34e == _io_insn_T[9:0] ? 32'h13 : _GEN_846; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_848 = 10'h34f == _io_insn_T[9:0] ? 32'h13 : _GEN_847; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_849 = 10'h350 == _io_insn_T[9:0] ? 32'h13 : _GEN_848; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_850 = 10'h351 == _io_insn_T[9:0] ? 32'h13 : _GEN_849; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_851 = 10'h352 == _io_insn_T[9:0] ? 32'h13 : _GEN_850; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_852 = 10'h353 == _io_insn_T[9:0] ? 32'h13 : _GEN_851; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_853 = 10'h354 == _io_insn_T[9:0] ? 32'h13 : _GEN_852; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_854 = 10'h355 == _io_insn_T[9:0] ? 32'h13 : _GEN_853; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_855 = 10'h356 == _io_insn_T[9:0] ? 32'h13 : _GEN_854; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_856 = 10'h357 == _io_insn_T[9:0] ? 32'h13 : _GEN_855; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_857 = 10'h358 == _io_insn_T[9:0] ? 32'h13 : _GEN_856; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_858 = 10'h359 == _io_insn_T[9:0] ? 32'h13 : _GEN_857; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_859 = 10'h35a == _io_insn_T[9:0] ? 32'h13 : _GEN_858; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_860 = 10'h35b == _io_insn_T[9:0] ? 32'h13 : _GEN_859; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_861 = 10'h35c == _io_insn_T[9:0] ? 32'h13 : _GEN_860; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_862 = 10'h35d == _io_insn_T[9:0] ? 32'h13 : _GEN_861; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_863 = 10'h35e == _io_insn_T[9:0] ? 32'h13 : _GEN_862; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_864 = 10'h35f == _io_insn_T[9:0] ? 32'h13 : _GEN_863; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_865 = 10'h360 == _io_insn_T[9:0] ? 32'h13 : _GEN_864; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_866 = 10'h361 == _io_insn_T[9:0] ? 32'h13 : _GEN_865; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_867 = 10'h362 == _io_insn_T[9:0] ? 32'h13 : _GEN_866; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_868 = 10'h363 == _io_insn_T[9:0] ? 32'h13 : _GEN_867; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_869 = 10'h364 == _io_insn_T[9:0] ? 32'h13 : _GEN_868; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_870 = 10'h365 == _io_insn_T[9:0] ? 32'h13 : _GEN_869; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_871 = 10'h366 == _io_insn_T[9:0] ? 32'h13 : _GEN_870; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_872 = 10'h367 == _io_insn_T[9:0] ? 32'h13 : _GEN_871; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_873 = 10'h368 == _io_insn_T[9:0] ? 32'h13 : _GEN_872; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_874 = 10'h369 == _io_insn_T[9:0] ? 32'h13 : _GEN_873; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_875 = 10'h36a == _io_insn_T[9:0] ? 32'h13 : _GEN_874; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_876 = 10'h36b == _io_insn_T[9:0] ? 32'h13 : _GEN_875; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_877 = 10'h36c == _io_insn_T[9:0] ? 32'h13 : _GEN_876; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_878 = 10'h36d == _io_insn_T[9:0] ? 32'h13 : _GEN_877; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_879 = 10'h36e == _io_insn_T[9:0] ? 32'h13 : _GEN_878; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_880 = 10'h36f == _io_insn_T[9:0] ? 32'h13 : _GEN_879; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_881 = 10'h370 == _io_insn_T[9:0] ? 32'h13 : _GEN_880; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_882 = 10'h371 == _io_insn_T[9:0] ? 32'h13 : _GEN_881; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_883 = 10'h372 == _io_insn_T[9:0] ? 32'h13 : _GEN_882; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_884 = 10'h373 == _io_insn_T[9:0] ? 32'h13 : _GEN_883; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_885 = 10'h374 == _io_insn_T[9:0] ? 32'h13 : _GEN_884; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_886 = 10'h375 == _io_insn_T[9:0] ? 32'h13 : _GEN_885; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_887 = 10'h376 == _io_insn_T[9:0] ? 32'h13 : _GEN_886; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_888 = 10'h377 == _io_insn_T[9:0] ? 32'h13 : _GEN_887; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_889 = 10'h378 == _io_insn_T[9:0] ? 32'h13 : _GEN_888; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_890 = 10'h379 == _io_insn_T[9:0] ? 32'h13 : _GEN_889; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_891 = 10'h37a == _io_insn_T[9:0] ? 32'h13 : _GEN_890; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_892 = 10'h37b == _io_insn_T[9:0] ? 32'h13 : _GEN_891; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_893 = 10'h37c == _io_insn_T[9:0] ? 32'h13 : _GEN_892; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_894 = 10'h37d == _io_insn_T[9:0] ? 32'h13 : _GEN_893; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_895 = 10'h37e == _io_insn_T[9:0] ? 32'h13 : _GEN_894; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_896 = 10'h37f == _io_insn_T[9:0] ? 32'h13 : _GEN_895; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_897 = 10'h380 == _io_insn_T[9:0] ? 32'h13 : _GEN_896; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_898 = 10'h381 == _io_insn_T[9:0] ? 32'h13 : _GEN_897; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_899 = 10'h382 == _io_insn_T[9:0] ? 32'h13 : _GEN_898; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_900 = 10'h383 == _io_insn_T[9:0] ? 32'h13 : _GEN_899; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_901 = 10'h384 == _io_insn_T[9:0] ? 32'h13 : _GEN_900; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_902 = 10'h385 == _io_insn_T[9:0] ? 32'h13 : _GEN_901; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_903 = 10'h386 == _io_insn_T[9:0] ? 32'h13 : _GEN_902; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_904 = 10'h387 == _io_insn_T[9:0] ? 32'h13 : _GEN_903; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_905 = 10'h388 == _io_insn_T[9:0] ? 32'h13 : _GEN_904; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_906 = 10'h389 == _io_insn_T[9:0] ? 32'h13 : _GEN_905; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_907 = 10'h38a == _io_insn_T[9:0] ? 32'h13 : _GEN_906; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_908 = 10'h38b == _io_insn_T[9:0] ? 32'h13 : _GEN_907; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_909 = 10'h38c == _io_insn_T[9:0] ? 32'h13 : _GEN_908; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_910 = 10'h38d == _io_insn_T[9:0] ? 32'h13 : _GEN_909; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_911 = 10'h38e == _io_insn_T[9:0] ? 32'h13 : _GEN_910; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_912 = 10'h38f == _io_insn_T[9:0] ? 32'h13 : _GEN_911; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_913 = 10'h390 == _io_insn_T[9:0] ? 32'h13 : _GEN_912; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_914 = 10'h391 == _io_insn_T[9:0] ? 32'h13 : _GEN_913; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_915 = 10'h392 == _io_insn_T[9:0] ? 32'h13 : _GEN_914; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_916 = 10'h393 == _io_insn_T[9:0] ? 32'h13 : _GEN_915; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_917 = 10'h394 == _io_insn_T[9:0] ? 32'h13 : _GEN_916; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_918 = 10'h395 == _io_insn_T[9:0] ? 32'h13 : _GEN_917; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_919 = 10'h396 == _io_insn_T[9:0] ? 32'h13 : _GEN_918; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_920 = 10'h397 == _io_insn_T[9:0] ? 32'h13 : _GEN_919; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_921 = 10'h398 == _io_insn_T[9:0] ? 32'h13 : _GEN_920; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_922 = 10'h399 == _io_insn_T[9:0] ? 32'h13 : _GEN_921; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_923 = 10'h39a == _io_insn_T[9:0] ? 32'h13 : _GEN_922; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_924 = 10'h39b == _io_insn_T[9:0] ? 32'h13 : _GEN_923; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_925 = 10'h39c == _io_insn_T[9:0] ? 32'h13 : _GEN_924; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_926 = 10'h39d == _io_insn_T[9:0] ? 32'h13 : _GEN_925; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_927 = 10'h39e == _io_insn_T[9:0] ? 32'h13 : _GEN_926; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_928 = 10'h39f == _io_insn_T[9:0] ? 32'h13 : _GEN_927; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_929 = 10'h3a0 == _io_insn_T[9:0] ? 32'h13 : _GEN_928; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_930 = 10'h3a1 == _io_insn_T[9:0] ? 32'h13 : _GEN_929; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_931 = 10'h3a2 == _io_insn_T[9:0] ? 32'h13 : _GEN_930; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_932 = 10'h3a3 == _io_insn_T[9:0] ? 32'h13 : _GEN_931; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_933 = 10'h3a4 == _io_insn_T[9:0] ? 32'h13 : _GEN_932; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_934 = 10'h3a5 == _io_insn_T[9:0] ? 32'h13 : _GEN_933; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_935 = 10'h3a6 == _io_insn_T[9:0] ? 32'h13 : _GEN_934; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_936 = 10'h3a7 == _io_insn_T[9:0] ? 32'h13 : _GEN_935; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_937 = 10'h3a8 == _io_insn_T[9:0] ? 32'h13 : _GEN_936; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_938 = 10'h3a9 == _io_insn_T[9:0] ? 32'h13 : _GEN_937; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_939 = 10'h3aa == _io_insn_T[9:0] ? 32'h13 : _GEN_938; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_940 = 10'h3ab == _io_insn_T[9:0] ? 32'h13 : _GEN_939; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_941 = 10'h3ac == _io_insn_T[9:0] ? 32'h13 : _GEN_940; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_942 = 10'h3ad == _io_insn_T[9:0] ? 32'h13 : _GEN_941; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_943 = 10'h3ae == _io_insn_T[9:0] ? 32'h13 : _GEN_942; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_944 = 10'h3af == _io_insn_T[9:0] ? 32'h13 : _GEN_943; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_945 = 10'h3b0 == _io_insn_T[9:0] ? 32'h13 : _GEN_944; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_946 = 10'h3b1 == _io_insn_T[9:0] ? 32'h13 : _GEN_945; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_947 = 10'h3b2 == _io_insn_T[9:0] ? 32'h13 : _GEN_946; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_948 = 10'h3b3 == _io_insn_T[9:0] ? 32'h13 : _GEN_947; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_949 = 10'h3b4 == _io_insn_T[9:0] ? 32'h13 : _GEN_948; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_950 = 10'h3b5 == _io_insn_T[9:0] ? 32'h13 : _GEN_949; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_951 = 10'h3b6 == _io_insn_T[9:0] ? 32'h13 : _GEN_950; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_952 = 10'h3b7 == _io_insn_T[9:0] ? 32'h13 : _GEN_951; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_953 = 10'h3b8 == _io_insn_T[9:0] ? 32'h13 : _GEN_952; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_954 = 10'h3b9 == _io_insn_T[9:0] ? 32'h13 : _GEN_953; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_955 = 10'h3ba == _io_insn_T[9:0] ? 32'h13 : _GEN_954; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_956 = 10'h3bb == _io_insn_T[9:0] ? 32'h13 : _GEN_955; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_957 = 10'h3bc == _io_insn_T[9:0] ? 32'h13 : _GEN_956; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_958 = 10'h3bd == _io_insn_T[9:0] ? 32'h13 : _GEN_957; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_959 = 10'h3be == _io_insn_T[9:0] ? 32'h13 : _GEN_958; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_960 = 10'h3bf == _io_insn_T[9:0] ? 32'h13 : _GEN_959; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_961 = 10'h3c0 == _io_insn_T[9:0] ? 32'h13 : _GEN_960; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_962 = 10'h3c1 == _io_insn_T[9:0] ? 32'h13 : _GEN_961; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_963 = 10'h3c2 == _io_insn_T[9:0] ? 32'h13 : _GEN_962; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_964 = 10'h3c3 == _io_insn_T[9:0] ? 32'h13 : _GEN_963; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_965 = 10'h3c4 == _io_insn_T[9:0] ? 32'h13 : _GEN_964; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_966 = 10'h3c5 == _io_insn_T[9:0] ? 32'h13 : _GEN_965; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_967 = 10'h3c6 == _io_insn_T[9:0] ? 32'h13 : _GEN_966; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_968 = 10'h3c7 == _io_insn_T[9:0] ? 32'h13 : _GEN_967; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_969 = 10'h3c8 == _io_insn_T[9:0] ? 32'h13 : _GEN_968; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_970 = 10'h3c9 == _io_insn_T[9:0] ? 32'h13 : _GEN_969; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_971 = 10'h3ca == _io_insn_T[9:0] ? 32'h13 : _GEN_970; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_972 = 10'h3cb == _io_insn_T[9:0] ? 32'h13 : _GEN_971; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_973 = 10'h3cc == _io_insn_T[9:0] ? 32'h13 : _GEN_972; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_974 = 10'h3cd == _io_insn_T[9:0] ? 32'h13 : _GEN_973; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_975 = 10'h3ce == _io_insn_T[9:0] ? 32'h13 : _GEN_974; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_976 = 10'h3cf == _io_insn_T[9:0] ? 32'h13 : _GEN_975; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_977 = 10'h3d0 == _io_insn_T[9:0] ? 32'h13 : _GEN_976; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_978 = 10'h3d1 == _io_insn_T[9:0] ? 32'h13 : _GEN_977; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_979 = 10'h3d2 == _io_insn_T[9:0] ? 32'h13 : _GEN_978; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_980 = 10'h3d3 == _io_insn_T[9:0] ? 32'h13 : _GEN_979; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_981 = 10'h3d4 == _io_insn_T[9:0] ? 32'h13 : _GEN_980; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_982 = 10'h3d5 == _io_insn_T[9:0] ? 32'h13 : _GEN_981; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_983 = 10'h3d6 == _io_insn_T[9:0] ? 32'h13 : _GEN_982; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_984 = 10'h3d7 == _io_insn_T[9:0] ? 32'h13 : _GEN_983; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_985 = 10'h3d8 == _io_insn_T[9:0] ? 32'h13 : _GEN_984; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_986 = 10'h3d9 == _io_insn_T[9:0] ? 32'h13 : _GEN_985; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_987 = 10'h3da == _io_insn_T[9:0] ? 32'h13 : _GEN_986; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_988 = 10'h3db == _io_insn_T[9:0] ? 32'h13 : _GEN_987; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_989 = 10'h3dc == _io_insn_T[9:0] ? 32'h13 : _GEN_988; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_990 = 10'h3dd == _io_insn_T[9:0] ? 32'h13 : _GEN_989; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_991 = 10'h3de == _io_insn_T[9:0] ? 32'h13 : _GEN_990; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_992 = 10'h3df == _io_insn_T[9:0] ? 32'h13 : _GEN_991; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_993 = 10'h3e0 == _io_insn_T[9:0] ? 32'h13 : _GEN_992; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_994 = 10'h3e1 == _io_insn_T[9:0] ? 32'h13 : _GEN_993; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_995 = 10'h3e2 == _io_insn_T[9:0] ? 32'h13 : _GEN_994; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_996 = 10'h3e3 == _io_insn_T[9:0] ? 32'h13 : _GEN_995; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_997 = 10'h3e4 == _io_insn_T[9:0] ? 32'h13 : _GEN_996; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_998 = 10'h3e5 == _io_insn_T[9:0] ? 32'h13 : _GEN_997; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_999 = 10'h3e6 == _io_insn_T[9:0] ? 32'h13 : _GEN_998; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1000 = 10'h3e7 == _io_insn_T[9:0] ? 32'h13 : _GEN_999; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1001 = 10'h3e8 == _io_insn_T[9:0] ? 32'h13 : _GEN_1000; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1002 = 10'h3e9 == _io_insn_T[9:0] ? 32'h13 : _GEN_1001; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1003 = 10'h3ea == _io_insn_T[9:0] ? 32'h13 : _GEN_1002; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1004 = 10'h3eb == _io_insn_T[9:0] ? 32'h13 : _GEN_1003; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1005 = 10'h3ec == _io_insn_T[9:0] ? 32'h13 : _GEN_1004; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1006 = 10'h3ed == _io_insn_T[9:0] ? 32'h13 : _GEN_1005; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1007 = 10'h3ee == _io_insn_T[9:0] ? 32'h13 : _GEN_1006; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1008 = 10'h3ef == _io_insn_T[9:0] ? 32'h13 : _GEN_1007; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1009 = 10'h3f0 == _io_insn_T[9:0] ? 32'h13 : _GEN_1008; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1010 = 10'h3f1 == _io_insn_T[9:0] ? 32'h13 : _GEN_1009; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1011 = 10'h3f2 == _io_insn_T[9:0] ? 32'h13 : _GEN_1010; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1012 = 10'h3f3 == _io_insn_T[9:0] ? 32'h13 : _GEN_1011; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1013 = 10'h3f4 == _io_insn_T[9:0] ? 32'h13 : _GEN_1012; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1014 = 10'h3f5 == _io_insn_T[9:0] ? 32'h13 : _GEN_1013; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1015 = 10'h3f6 == _io_insn_T[9:0] ? 32'h13 : _GEN_1014; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1016 = 10'h3f7 == _io_insn_T[9:0] ? 32'h13 : _GEN_1015; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1017 = 10'h3f8 == _io_insn_T[9:0] ? 32'h13 : _GEN_1016; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1018 = 10'h3f9 == _io_insn_T[9:0] ? 32'h13 : _GEN_1017; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1019 = 10'h3fa == _io_insn_T[9:0] ? 32'h13 : _GEN_1018; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1020 = 10'h3fb == _io_insn_T[9:0] ? 32'h13 : _GEN_1019; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1021 = 10'h3fc == _io_insn_T[9:0] ? 32'h13 : _GEN_1020; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1022 = 10'h3fd == _io_insn_T[9:0] ? 32'h13 : _GEN_1021; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1023 = 10'h3fe == _io_insn_T[9:0] ? 32'h13 : _GEN_1022; // @[cpu.scala 45:{13,13}]
  wire [31:0] _GEN_1024 = 10'h3ff == _io_insn_T[9:0] ? 32'h13 : _GEN_1023; // @[cpu.scala 45:{13,13}]
  assign io_nPC = counterReg == 2'h1 ? _io_nPC_T_1 : io_PC; // @[cpu.scala 43:26 44:12 47:12]
  assign io_insn = counterReg == 2'h1 ? _GEN_1024 : 32'h13; // @[cpu.scala 43:26 45:13 48:13]
  always @(posedge clock) begin
    if (reset) begin // @[cpu.scala 37:27]
      counterReg <= 2'h0; // @[cpu.scala 37:27]
    end else if (io_reset) begin // @[cpu.scala 38:18]
      counterReg <= 2'h0; // @[cpu.scala 39:16]
    end else begin
      counterReg <= _counterReg_T_1; // @[cpu.scala 41:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counterReg = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RISCVCPUv2Bubble(
  input         clock,
  input         reset,
  input         io_rvfi_rst,
  input  [31:0] io_rvfi_insn_in_0,
  input  [31:0] io_rvfi_insn_in_1,
  output [63:0] io_rvfi_regs_0,
  output [63:0] io_rvfi_regs_1,
  output [63:0] io_rvfi_regs_2,
  output [63:0] io_rvfi_regs_3,
  output [63:0] io_rvfi_regs_4,
  output [63:0] io_rvfi_regs_5,
  output [63:0] io_rvfi_regs_6,
  output [63:0] io_rvfi_regs_7,
  output [63:0] io_rvfi_regs_8,
  output [63:0] io_rvfi_regs_9,
  output [63:0] io_rvfi_regs_10,
  output [63:0] io_rvfi_regs_11,
  output [63:0] io_rvfi_regs_12,
  output [63:0] io_rvfi_regs_13,
  output [63:0] io_rvfi_regs_14,
  output [63:0] io_rvfi_regs_15,
  output [63:0] io_rvfi_regs_16,
  output [63:0] io_rvfi_regs_17,
  output [63:0] io_rvfi_regs_18,
  output [63:0] io_rvfi_regs_19,
  output [63:0] io_rvfi_regs_20,
  output [63:0] io_rvfi_regs_21,
  output [63:0] io_rvfi_regs_22,
  output [63:0] io_rvfi_regs_23,
  output [63:0] io_rvfi_regs_24,
  output [63:0] io_rvfi_regs_25,
  output [63:0] io_rvfi_regs_26,
  output [63:0] io_rvfi_regs_27,
  output [63:0] io_rvfi_regs_28,
  output [63:0] io_rvfi_regs_29,
  output [63:0] io_rvfi_regs_30,
  output [63:0] io_rvfi_regs_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [63:0] _RAND_1068;
`endif // RANDOMIZE_REG_INIT
  wire  ControlUnit_clock; // @[cpu.scala 293:20]
  wire  ControlUnit_reset; // @[cpu.scala 293:20]
  wire  ControlUnit_io_reset; // @[cpu.scala 293:20]
  wire [31:0] ControlUnit_io_insns_0; // @[cpu.scala 293:20]
  wire [31:0] ControlUnit_io_insns_1; // @[cpu.scala 293:20]
  wire [63:0] ControlUnit_io_PC; // @[cpu.scala 293:20]
  wire [63:0] ControlUnit_io_nPC; // @[cpu.scala 293:20]
  wire [31:0] ControlUnit_io_insn; // @[cpu.scala 293:20]
  reg [63:0] PC; // @[cpu.scala 277:19]
  reg [63:0] Regs_0; // @[cpu.scala 278:21]
  reg [63:0] Regs_1; // @[cpu.scala 278:21]
  reg [63:0] Regs_2; // @[cpu.scala 278:21]
  reg [63:0] Regs_3; // @[cpu.scala 278:21]
  reg [63:0] Regs_4; // @[cpu.scala 278:21]
  reg [63:0] Regs_5; // @[cpu.scala 278:21]
  reg [63:0] Regs_6; // @[cpu.scala 278:21]
  reg [63:0] Regs_7; // @[cpu.scala 278:21]
  reg [63:0] Regs_8; // @[cpu.scala 278:21]
  reg [63:0] Regs_9; // @[cpu.scala 278:21]
  reg [63:0] Regs_10; // @[cpu.scala 278:21]
  reg [63:0] Regs_11; // @[cpu.scala 278:21]
  reg [63:0] Regs_12; // @[cpu.scala 278:21]
  reg [63:0] Regs_13; // @[cpu.scala 278:21]
  reg [63:0] Regs_14; // @[cpu.scala 278:21]
  reg [63:0] Regs_15; // @[cpu.scala 278:21]
  reg [63:0] Regs_16; // @[cpu.scala 278:21]
  reg [63:0] Regs_17; // @[cpu.scala 278:21]
  reg [63:0] Regs_18; // @[cpu.scala 278:21]
  reg [63:0] Regs_19; // @[cpu.scala 278:21]
  reg [63:0] Regs_20; // @[cpu.scala 278:21]
  reg [63:0] Regs_21; // @[cpu.scala 278:21]
  reg [63:0] Regs_22; // @[cpu.scala 278:21]
  reg [63:0] Regs_23; // @[cpu.scala 278:21]
  reg [63:0] Regs_24; // @[cpu.scala 278:21]
  reg [63:0] Regs_25; // @[cpu.scala 278:21]
  reg [63:0] Regs_26; // @[cpu.scala 278:21]
  reg [63:0] Regs_27; // @[cpu.scala 278:21]
  reg [63:0] Regs_28; // @[cpu.scala 278:21]
  reg [63:0] Regs_29; // @[cpu.scala 278:21]
  reg [63:0] Regs_30; // @[cpu.scala 278:21]
  reg [63:0] Regs_31; // @[cpu.scala 278:21]
  reg [63:0] IDEXA; // @[cpu.scala 280:58]
  reg [63:0] IDEXB; // @[cpu.scala 280:58]
  reg [63:0] EXMEMB; // @[cpu.scala 280:58]
  reg [63:0] EXMEMALUOut; // @[cpu.scala 280:58]
  reg [63:0] MEMWBValue; // @[cpu.scala 280:58]
  reg [31:0] DMemory_0; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1; // @[cpu.scala 282:24]
  reg [31:0] DMemory_2; // @[cpu.scala 282:24]
  reg [31:0] DMemory_3; // @[cpu.scala 282:24]
  reg [31:0] DMemory_4; // @[cpu.scala 282:24]
  reg [31:0] DMemory_5; // @[cpu.scala 282:24]
  reg [31:0] DMemory_6; // @[cpu.scala 282:24]
  reg [31:0] DMemory_7; // @[cpu.scala 282:24]
  reg [31:0] DMemory_8; // @[cpu.scala 282:24]
  reg [31:0] DMemory_9; // @[cpu.scala 282:24]
  reg [31:0] DMemory_10; // @[cpu.scala 282:24]
  reg [31:0] DMemory_11; // @[cpu.scala 282:24]
  reg [31:0] DMemory_12; // @[cpu.scala 282:24]
  reg [31:0] DMemory_13; // @[cpu.scala 282:24]
  reg [31:0] DMemory_14; // @[cpu.scala 282:24]
  reg [31:0] DMemory_15; // @[cpu.scala 282:24]
  reg [31:0] DMemory_16; // @[cpu.scala 282:24]
  reg [31:0] DMemory_17; // @[cpu.scala 282:24]
  reg [31:0] DMemory_18; // @[cpu.scala 282:24]
  reg [31:0] DMemory_19; // @[cpu.scala 282:24]
  reg [31:0] DMemory_20; // @[cpu.scala 282:24]
  reg [31:0] DMemory_21; // @[cpu.scala 282:24]
  reg [31:0] DMemory_22; // @[cpu.scala 282:24]
  reg [31:0] DMemory_23; // @[cpu.scala 282:24]
  reg [31:0] DMemory_24; // @[cpu.scala 282:24]
  reg [31:0] DMemory_25; // @[cpu.scala 282:24]
  reg [31:0] DMemory_26; // @[cpu.scala 282:24]
  reg [31:0] DMemory_27; // @[cpu.scala 282:24]
  reg [31:0] DMemory_28; // @[cpu.scala 282:24]
  reg [31:0] DMemory_29; // @[cpu.scala 282:24]
  reg [31:0] DMemory_30; // @[cpu.scala 282:24]
  reg [31:0] DMemory_31; // @[cpu.scala 282:24]
  reg [31:0] DMemory_32; // @[cpu.scala 282:24]
  reg [31:0] DMemory_33; // @[cpu.scala 282:24]
  reg [31:0] DMemory_34; // @[cpu.scala 282:24]
  reg [31:0] DMemory_35; // @[cpu.scala 282:24]
  reg [31:0] DMemory_36; // @[cpu.scala 282:24]
  reg [31:0] DMemory_37; // @[cpu.scala 282:24]
  reg [31:0] DMemory_38; // @[cpu.scala 282:24]
  reg [31:0] DMemory_39; // @[cpu.scala 282:24]
  reg [31:0] DMemory_40; // @[cpu.scala 282:24]
  reg [31:0] DMemory_41; // @[cpu.scala 282:24]
  reg [31:0] DMemory_42; // @[cpu.scala 282:24]
  reg [31:0] DMemory_43; // @[cpu.scala 282:24]
  reg [31:0] DMemory_44; // @[cpu.scala 282:24]
  reg [31:0] DMemory_45; // @[cpu.scala 282:24]
  reg [31:0] DMemory_46; // @[cpu.scala 282:24]
  reg [31:0] DMemory_47; // @[cpu.scala 282:24]
  reg [31:0] DMemory_48; // @[cpu.scala 282:24]
  reg [31:0] DMemory_49; // @[cpu.scala 282:24]
  reg [31:0] DMemory_50; // @[cpu.scala 282:24]
  reg [31:0] DMemory_51; // @[cpu.scala 282:24]
  reg [31:0] DMemory_52; // @[cpu.scala 282:24]
  reg [31:0] DMemory_53; // @[cpu.scala 282:24]
  reg [31:0] DMemory_54; // @[cpu.scala 282:24]
  reg [31:0] DMemory_55; // @[cpu.scala 282:24]
  reg [31:0] DMemory_56; // @[cpu.scala 282:24]
  reg [31:0] DMemory_57; // @[cpu.scala 282:24]
  reg [31:0] DMemory_58; // @[cpu.scala 282:24]
  reg [31:0] DMemory_59; // @[cpu.scala 282:24]
  reg [31:0] DMemory_60; // @[cpu.scala 282:24]
  reg [31:0] DMemory_61; // @[cpu.scala 282:24]
  reg [31:0] DMemory_62; // @[cpu.scala 282:24]
  reg [31:0] DMemory_63; // @[cpu.scala 282:24]
  reg [31:0] DMemory_64; // @[cpu.scala 282:24]
  reg [31:0] DMemory_65; // @[cpu.scala 282:24]
  reg [31:0] DMemory_66; // @[cpu.scala 282:24]
  reg [31:0] DMemory_67; // @[cpu.scala 282:24]
  reg [31:0] DMemory_68; // @[cpu.scala 282:24]
  reg [31:0] DMemory_69; // @[cpu.scala 282:24]
  reg [31:0] DMemory_70; // @[cpu.scala 282:24]
  reg [31:0] DMemory_71; // @[cpu.scala 282:24]
  reg [31:0] DMemory_72; // @[cpu.scala 282:24]
  reg [31:0] DMemory_73; // @[cpu.scala 282:24]
  reg [31:0] DMemory_74; // @[cpu.scala 282:24]
  reg [31:0] DMemory_75; // @[cpu.scala 282:24]
  reg [31:0] DMemory_76; // @[cpu.scala 282:24]
  reg [31:0] DMemory_77; // @[cpu.scala 282:24]
  reg [31:0] DMemory_78; // @[cpu.scala 282:24]
  reg [31:0] DMemory_79; // @[cpu.scala 282:24]
  reg [31:0] DMemory_80; // @[cpu.scala 282:24]
  reg [31:0] DMemory_81; // @[cpu.scala 282:24]
  reg [31:0] DMemory_82; // @[cpu.scala 282:24]
  reg [31:0] DMemory_83; // @[cpu.scala 282:24]
  reg [31:0] DMemory_84; // @[cpu.scala 282:24]
  reg [31:0] DMemory_85; // @[cpu.scala 282:24]
  reg [31:0] DMemory_86; // @[cpu.scala 282:24]
  reg [31:0] DMemory_87; // @[cpu.scala 282:24]
  reg [31:0] DMemory_88; // @[cpu.scala 282:24]
  reg [31:0] DMemory_89; // @[cpu.scala 282:24]
  reg [31:0] DMemory_90; // @[cpu.scala 282:24]
  reg [31:0] DMemory_91; // @[cpu.scala 282:24]
  reg [31:0] DMemory_92; // @[cpu.scala 282:24]
  reg [31:0] DMemory_93; // @[cpu.scala 282:24]
  reg [31:0] DMemory_94; // @[cpu.scala 282:24]
  reg [31:0] DMemory_95; // @[cpu.scala 282:24]
  reg [31:0] DMemory_96; // @[cpu.scala 282:24]
  reg [31:0] DMemory_97; // @[cpu.scala 282:24]
  reg [31:0] DMemory_98; // @[cpu.scala 282:24]
  reg [31:0] DMemory_99; // @[cpu.scala 282:24]
  reg [31:0] DMemory_100; // @[cpu.scala 282:24]
  reg [31:0] DMemory_101; // @[cpu.scala 282:24]
  reg [31:0] DMemory_102; // @[cpu.scala 282:24]
  reg [31:0] DMemory_103; // @[cpu.scala 282:24]
  reg [31:0] DMemory_104; // @[cpu.scala 282:24]
  reg [31:0] DMemory_105; // @[cpu.scala 282:24]
  reg [31:0] DMemory_106; // @[cpu.scala 282:24]
  reg [31:0] DMemory_107; // @[cpu.scala 282:24]
  reg [31:0] DMemory_108; // @[cpu.scala 282:24]
  reg [31:0] DMemory_109; // @[cpu.scala 282:24]
  reg [31:0] DMemory_110; // @[cpu.scala 282:24]
  reg [31:0] DMemory_111; // @[cpu.scala 282:24]
  reg [31:0] DMemory_112; // @[cpu.scala 282:24]
  reg [31:0] DMemory_113; // @[cpu.scala 282:24]
  reg [31:0] DMemory_114; // @[cpu.scala 282:24]
  reg [31:0] DMemory_115; // @[cpu.scala 282:24]
  reg [31:0] DMemory_116; // @[cpu.scala 282:24]
  reg [31:0] DMemory_117; // @[cpu.scala 282:24]
  reg [31:0] DMemory_118; // @[cpu.scala 282:24]
  reg [31:0] DMemory_119; // @[cpu.scala 282:24]
  reg [31:0] DMemory_120; // @[cpu.scala 282:24]
  reg [31:0] DMemory_121; // @[cpu.scala 282:24]
  reg [31:0] DMemory_122; // @[cpu.scala 282:24]
  reg [31:0] DMemory_123; // @[cpu.scala 282:24]
  reg [31:0] DMemory_124; // @[cpu.scala 282:24]
  reg [31:0] DMemory_125; // @[cpu.scala 282:24]
  reg [31:0] DMemory_126; // @[cpu.scala 282:24]
  reg [31:0] DMemory_127; // @[cpu.scala 282:24]
  reg [31:0] DMemory_128; // @[cpu.scala 282:24]
  reg [31:0] DMemory_129; // @[cpu.scala 282:24]
  reg [31:0] DMemory_130; // @[cpu.scala 282:24]
  reg [31:0] DMemory_131; // @[cpu.scala 282:24]
  reg [31:0] DMemory_132; // @[cpu.scala 282:24]
  reg [31:0] DMemory_133; // @[cpu.scala 282:24]
  reg [31:0] DMemory_134; // @[cpu.scala 282:24]
  reg [31:0] DMemory_135; // @[cpu.scala 282:24]
  reg [31:0] DMemory_136; // @[cpu.scala 282:24]
  reg [31:0] DMemory_137; // @[cpu.scala 282:24]
  reg [31:0] DMemory_138; // @[cpu.scala 282:24]
  reg [31:0] DMemory_139; // @[cpu.scala 282:24]
  reg [31:0] DMemory_140; // @[cpu.scala 282:24]
  reg [31:0] DMemory_141; // @[cpu.scala 282:24]
  reg [31:0] DMemory_142; // @[cpu.scala 282:24]
  reg [31:0] DMemory_143; // @[cpu.scala 282:24]
  reg [31:0] DMemory_144; // @[cpu.scala 282:24]
  reg [31:0] DMemory_145; // @[cpu.scala 282:24]
  reg [31:0] DMemory_146; // @[cpu.scala 282:24]
  reg [31:0] DMemory_147; // @[cpu.scala 282:24]
  reg [31:0] DMemory_148; // @[cpu.scala 282:24]
  reg [31:0] DMemory_149; // @[cpu.scala 282:24]
  reg [31:0] DMemory_150; // @[cpu.scala 282:24]
  reg [31:0] DMemory_151; // @[cpu.scala 282:24]
  reg [31:0] DMemory_152; // @[cpu.scala 282:24]
  reg [31:0] DMemory_153; // @[cpu.scala 282:24]
  reg [31:0] DMemory_154; // @[cpu.scala 282:24]
  reg [31:0] DMemory_155; // @[cpu.scala 282:24]
  reg [31:0] DMemory_156; // @[cpu.scala 282:24]
  reg [31:0] DMemory_157; // @[cpu.scala 282:24]
  reg [31:0] DMemory_158; // @[cpu.scala 282:24]
  reg [31:0] DMemory_159; // @[cpu.scala 282:24]
  reg [31:0] DMemory_160; // @[cpu.scala 282:24]
  reg [31:0] DMemory_161; // @[cpu.scala 282:24]
  reg [31:0] DMemory_162; // @[cpu.scala 282:24]
  reg [31:0] DMemory_163; // @[cpu.scala 282:24]
  reg [31:0] DMemory_164; // @[cpu.scala 282:24]
  reg [31:0] DMemory_165; // @[cpu.scala 282:24]
  reg [31:0] DMemory_166; // @[cpu.scala 282:24]
  reg [31:0] DMemory_167; // @[cpu.scala 282:24]
  reg [31:0] DMemory_168; // @[cpu.scala 282:24]
  reg [31:0] DMemory_169; // @[cpu.scala 282:24]
  reg [31:0] DMemory_170; // @[cpu.scala 282:24]
  reg [31:0] DMemory_171; // @[cpu.scala 282:24]
  reg [31:0] DMemory_172; // @[cpu.scala 282:24]
  reg [31:0] DMemory_173; // @[cpu.scala 282:24]
  reg [31:0] DMemory_174; // @[cpu.scala 282:24]
  reg [31:0] DMemory_175; // @[cpu.scala 282:24]
  reg [31:0] DMemory_176; // @[cpu.scala 282:24]
  reg [31:0] DMemory_177; // @[cpu.scala 282:24]
  reg [31:0] DMemory_178; // @[cpu.scala 282:24]
  reg [31:0] DMemory_179; // @[cpu.scala 282:24]
  reg [31:0] DMemory_180; // @[cpu.scala 282:24]
  reg [31:0] DMemory_181; // @[cpu.scala 282:24]
  reg [31:0] DMemory_182; // @[cpu.scala 282:24]
  reg [31:0] DMemory_183; // @[cpu.scala 282:24]
  reg [31:0] DMemory_184; // @[cpu.scala 282:24]
  reg [31:0] DMemory_185; // @[cpu.scala 282:24]
  reg [31:0] DMemory_186; // @[cpu.scala 282:24]
  reg [31:0] DMemory_187; // @[cpu.scala 282:24]
  reg [31:0] DMemory_188; // @[cpu.scala 282:24]
  reg [31:0] DMemory_189; // @[cpu.scala 282:24]
  reg [31:0] DMemory_190; // @[cpu.scala 282:24]
  reg [31:0] DMemory_191; // @[cpu.scala 282:24]
  reg [31:0] DMemory_192; // @[cpu.scala 282:24]
  reg [31:0] DMemory_193; // @[cpu.scala 282:24]
  reg [31:0] DMemory_194; // @[cpu.scala 282:24]
  reg [31:0] DMemory_195; // @[cpu.scala 282:24]
  reg [31:0] DMemory_196; // @[cpu.scala 282:24]
  reg [31:0] DMemory_197; // @[cpu.scala 282:24]
  reg [31:0] DMemory_198; // @[cpu.scala 282:24]
  reg [31:0] DMemory_199; // @[cpu.scala 282:24]
  reg [31:0] DMemory_200; // @[cpu.scala 282:24]
  reg [31:0] DMemory_201; // @[cpu.scala 282:24]
  reg [31:0] DMemory_202; // @[cpu.scala 282:24]
  reg [31:0] DMemory_203; // @[cpu.scala 282:24]
  reg [31:0] DMemory_204; // @[cpu.scala 282:24]
  reg [31:0] DMemory_205; // @[cpu.scala 282:24]
  reg [31:0] DMemory_206; // @[cpu.scala 282:24]
  reg [31:0] DMemory_207; // @[cpu.scala 282:24]
  reg [31:0] DMemory_208; // @[cpu.scala 282:24]
  reg [31:0] DMemory_209; // @[cpu.scala 282:24]
  reg [31:0] DMemory_210; // @[cpu.scala 282:24]
  reg [31:0] DMemory_211; // @[cpu.scala 282:24]
  reg [31:0] DMemory_212; // @[cpu.scala 282:24]
  reg [31:0] DMemory_213; // @[cpu.scala 282:24]
  reg [31:0] DMemory_214; // @[cpu.scala 282:24]
  reg [31:0] DMemory_215; // @[cpu.scala 282:24]
  reg [31:0] DMemory_216; // @[cpu.scala 282:24]
  reg [31:0] DMemory_217; // @[cpu.scala 282:24]
  reg [31:0] DMemory_218; // @[cpu.scala 282:24]
  reg [31:0] DMemory_219; // @[cpu.scala 282:24]
  reg [31:0] DMemory_220; // @[cpu.scala 282:24]
  reg [31:0] DMemory_221; // @[cpu.scala 282:24]
  reg [31:0] DMemory_222; // @[cpu.scala 282:24]
  reg [31:0] DMemory_223; // @[cpu.scala 282:24]
  reg [31:0] DMemory_224; // @[cpu.scala 282:24]
  reg [31:0] DMemory_225; // @[cpu.scala 282:24]
  reg [31:0] DMemory_226; // @[cpu.scala 282:24]
  reg [31:0] DMemory_227; // @[cpu.scala 282:24]
  reg [31:0] DMemory_228; // @[cpu.scala 282:24]
  reg [31:0] DMemory_229; // @[cpu.scala 282:24]
  reg [31:0] DMemory_230; // @[cpu.scala 282:24]
  reg [31:0] DMemory_231; // @[cpu.scala 282:24]
  reg [31:0] DMemory_232; // @[cpu.scala 282:24]
  reg [31:0] DMemory_233; // @[cpu.scala 282:24]
  reg [31:0] DMemory_234; // @[cpu.scala 282:24]
  reg [31:0] DMemory_235; // @[cpu.scala 282:24]
  reg [31:0] DMemory_236; // @[cpu.scala 282:24]
  reg [31:0] DMemory_237; // @[cpu.scala 282:24]
  reg [31:0] DMemory_238; // @[cpu.scala 282:24]
  reg [31:0] DMemory_239; // @[cpu.scala 282:24]
  reg [31:0] DMemory_240; // @[cpu.scala 282:24]
  reg [31:0] DMemory_241; // @[cpu.scala 282:24]
  reg [31:0] DMemory_242; // @[cpu.scala 282:24]
  reg [31:0] DMemory_243; // @[cpu.scala 282:24]
  reg [31:0] DMemory_244; // @[cpu.scala 282:24]
  reg [31:0] DMemory_245; // @[cpu.scala 282:24]
  reg [31:0] DMemory_246; // @[cpu.scala 282:24]
  reg [31:0] DMemory_247; // @[cpu.scala 282:24]
  reg [31:0] DMemory_248; // @[cpu.scala 282:24]
  reg [31:0] DMemory_249; // @[cpu.scala 282:24]
  reg [31:0] DMemory_250; // @[cpu.scala 282:24]
  reg [31:0] DMemory_251; // @[cpu.scala 282:24]
  reg [31:0] DMemory_252; // @[cpu.scala 282:24]
  reg [31:0] DMemory_253; // @[cpu.scala 282:24]
  reg [31:0] DMemory_254; // @[cpu.scala 282:24]
  reg [31:0] DMemory_255; // @[cpu.scala 282:24]
  reg [31:0] DMemory_256; // @[cpu.scala 282:24]
  reg [31:0] DMemory_257; // @[cpu.scala 282:24]
  reg [31:0] DMemory_258; // @[cpu.scala 282:24]
  reg [31:0] DMemory_259; // @[cpu.scala 282:24]
  reg [31:0] DMemory_260; // @[cpu.scala 282:24]
  reg [31:0] DMemory_261; // @[cpu.scala 282:24]
  reg [31:0] DMemory_262; // @[cpu.scala 282:24]
  reg [31:0] DMemory_263; // @[cpu.scala 282:24]
  reg [31:0] DMemory_264; // @[cpu.scala 282:24]
  reg [31:0] DMemory_265; // @[cpu.scala 282:24]
  reg [31:0] DMemory_266; // @[cpu.scala 282:24]
  reg [31:0] DMemory_267; // @[cpu.scala 282:24]
  reg [31:0] DMemory_268; // @[cpu.scala 282:24]
  reg [31:0] DMemory_269; // @[cpu.scala 282:24]
  reg [31:0] DMemory_270; // @[cpu.scala 282:24]
  reg [31:0] DMemory_271; // @[cpu.scala 282:24]
  reg [31:0] DMemory_272; // @[cpu.scala 282:24]
  reg [31:0] DMemory_273; // @[cpu.scala 282:24]
  reg [31:0] DMemory_274; // @[cpu.scala 282:24]
  reg [31:0] DMemory_275; // @[cpu.scala 282:24]
  reg [31:0] DMemory_276; // @[cpu.scala 282:24]
  reg [31:0] DMemory_277; // @[cpu.scala 282:24]
  reg [31:0] DMemory_278; // @[cpu.scala 282:24]
  reg [31:0] DMemory_279; // @[cpu.scala 282:24]
  reg [31:0] DMemory_280; // @[cpu.scala 282:24]
  reg [31:0] DMemory_281; // @[cpu.scala 282:24]
  reg [31:0] DMemory_282; // @[cpu.scala 282:24]
  reg [31:0] DMemory_283; // @[cpu.scala 282:24]
  reg [31:0] DMemory_284; // @[cpu.scala 282:24]
  reg [31:0] DMemory_285; // @[cpu.scala 282:24]
  reg [31:0] DMemory_286; // @[cpu.scala 282:24]
  reg [31:0] DMemory_287; // @[cpu.scala 282:24]
  reg [31:0] DMemory_288; // @[cpu.scala 282:24]
  reg [31:0] DMemory_289; // @[cpu.scala 282:24]
  reg [31:0] DMemory_290; // @[cpu.scala 282:24]
  reg [31:0] DMemory_291; // @[cpu.scala 282:24]
  reg [31:0] DMemory_292; // @[cpu.scala 282:24]
  reg [31:0] DMemory_293; // @[cpu.scala 282:24]
  reg [31:0] DMemory_294; // @[cpu.scala 282:24]
  reg [31:0] DMemory_295; // @[cpu.scala 282:24]
  reg [31:0] DMemory_296; // @[cpu.scala 282:24]
  reg [31:0] DMemory_297; // @[cpu.scala 282:24]
  reg [31:0] DMemory_298; // @[cpu.scala 282:24]
  reg [31:0] DMemory_299; // @[cpu.scala 282:24]
  reg [31:0] DMemory_300; // @[cpu.scala 282:24]
  reg [31:0] DMemory_301; // @[cpu.scala 282:24]
  reg [31:0] DMemory_302; // @[cpu.scala 282:24]
  reg [31:0] DMemory_303; // @[cpu.scala 282:24]
  reg [31:0] DMemory_304; // @[cpu.scala 282:24]
  reg [31:0] DMemory_305; // @[cpu.scala 282:24]
  reg [31:0] DMemory_306; // @[cpu.scala 282:24]
  reg [31:0] DMemory_307; // @[cpu.scala 282:24]
  reg [31:0] DMemory_308; // @[cpu.scala 282:24]
  reg [31:0] DMemory_309; // @[cpu.scala 282:24]
  reg [31:0] DMemory_310; // @[cpu.scala 282:24]
  reg [31:0] DMemory_311; // @[cpu.scala 282:24]
  reg [31:0] DMemory_312; // @[cpu.scala 282:24]
  reg [31:0] DMemory_313; // @[cpu.scala 282:24]
  reg [31:0] DMemory_314; // @[cpu.scala 282:24]
  reg [31:0] DMemory_315; // @[cpu.scala 282:24]
  reg [31:0] DMemory_316; // @[cpu.scala 282:24]
  reg [31:0] DMemory_317; // @[cpu.scala 282:24]
  reg [31:0] DMemory_318; // @[cpu.scala 282:24]
  reg [31:0] DMemory_319; // @[cpu.scala 282:24]
  reg [31:0] DMemory_320; // @[cpu.scala 282:24]
  reg [31:0] DMemory_321; // @[cpu.scala 282:24]
  reg [31:0] DMemory_322; // @[cpu.scala 282:24]
  reg [31:0] DMemory_323; // @[cpu.scala 282:24]
  reg [31:0] DMemory_324; // @[cpu.scala 282:24]
  reg [31:0] DMemory_325; // @[cpu.scala 282:24]
  reg [31:0] DMemory_326; // @[cpu.scala 282:24]
  reg [31:0] DMemory_327; // @[cpu.scala 282:24]
  reg [31:0] DMemory_328; // @[cpu.scala 282:24]
  reg [31:0] DMemory_329; // @[cpu.scala 282:24]
  reg [31:0] DMemory_330; // @[cpu.scala 282:24]
  reg [31:0] DMemory_331; // @[cpu.scala 282:24]
  reg [31:0] DMemory_332; // @[cpu.scala 282:24]
  reg [31:0] DMemory_333; // @[cpu.scala 282:24]
  reg [31:0] DMemory_334; // @[cpu.scala 282:24]
  reg [31:0] DMemory_335; // @[cpu.scala 282:24]
  reg [31:0] DMemory_336; // @[cpu.scala 282:24]
  reg [31:0] DMemory_337; // @[cpu.scala 282:24]
  reg [31:0] DMemory_338; // @[cpu.scala 282:24]
  reg [31:0] DMemory_339; // @[cpu.scala 282:24]
  reg [31:0] DMemory_340; // @[cpu.scala 282:24]
  reg [31:0] DMemory_341; // @[cpu.scala 282:24]
  reg [31:0] DMemory_342; // @[cpu.scala 282:24]
  reg [31:0] DMemory_343; // @[cpu.scala 282:24]
  reg [31:0] DMemory_344; // @[cpu.scala 282:24]
  reg [31:0] DMemory_345; // @[cpu.scala 282:24]
  reg [31:0] DMemory_346; // @[cpu.scala 282:24]
  reg [31:0] DMemory_347; // @[cpu.scala 282:24]
  reg [31:0] DMemory_348; // @[cpu.scala 282:24]
  reg [31:0] DMemory_349; // @[cpu.scala 282:24]
  reg [31:0] DMemory_350; // @[cpu.scala 282:24]
  reg [31:0] DMemory_351; // @[cpu.scala 282:24]
  reg [31:0] DMemory_352; // @[cpu.scala 282:24]
  reg [31:0] DMemory_353; // @[cpu.scala 282:24]
  reg [31:0] DMemory_354; // @[cpu.scala 282:24]
  reg [31:0] DMemory_355; // @[cpu.scala 282:24]
  reg [31:0] DMemory_356; // @[cpu.scala 282:24]
  reg [31:0] DMemory_357; // @[cpu.scala 282:24]
  reg [31:0] DMemory_358; // @[cpu.scala 282:24]
  reg [31:0] DMemory_359; // @[cpu.scala 282:24]
  reg [31:0] DMemory_360; // @[cpu.scala 282:24]
  reg [31:0] DMemory_361; // @[cpu.scala 282:24]
  reg [31:0] DMemory_362; // @[cpu.scala 282:24]
  reg [31:0] DMemory_363; // @[cpu.scala 282:24]
  reg [31:0] DMemory_364; // @[cpu.scala 282:24]
  reg [31:0] DMemory_365; // @[cpu.scala 282:24]
  reg [31:0] DMemory_366; // @[cpu.scala 282:24]
  reg [31:0] DMemory_367; // @[cpu.scala 282:24]
  reg [31:0] DMemory_368; // @[cpu.scala 282:24]
  reg [31:0] DMemory_369; // @[cpu.scala 282:24]
  reg [31:0] DMemory_370; // @[cpu.scala 282:24]
  reg [31:0] DMemory_371; // @[cpu.scala 282:24]
  reg [31:0] DMemory_372; // @[cpu.scala 282:24]
  reg [31:0] DMemory_373; // @[cpu.scala 282:24]
  reg [31:0] DMemory_374; // @[cpu.scala 282:24]
  reg [31:0] DMemory_375; // @[cpu.scala 282:24]
  reg [31:0] DMemory_376; // @[cpu.scala 282:24]
  reg [31:0] DMemory_377; // @[cpu.scala 282:24]
  reg [31:0] DMemory_378; // @[cpu.scala 282:24]
  reg [31:0] DMemory_379; // @[cpu.scala 282:24]
  reg [31:0] DMemory_380; // @[cpu.scala 282:24]
  reg [31:0] DMemory_381; // @[cpu.scala 282:24]
  reg [31:0] DMemory_382; // @[cpu.scala 282:24]
  reg [31:0] DMemory_383; // @[cpu.scala 282:24]
  reg [31:0] DMemory_384; // @[cpu.scala 282:24]
  reg [31:0] DMemory_385; // @[cpu.scala 282:24]
  reg [31:0] DMemory_386; // @[cpu.scala 282:24]
  reg [31:0] DMemory_387; // @[cpu.scala 282:24]
  reg [31:0] DMemory_388; // @[cpu.scala 282:24]
  reg [31:0] DMemory_389; // @[cpu.scala 282:24]
  reg [31:0] DMemory_390; // @[cpu.scala 282:24]
  reg [31:0] DMemory_391; // @[cpu.scala 282:24]
  reg [31:0] DMemory_392; // @[cpu.scala 282:24]
  reg [31:0] DMemory_393; // @[cpu.scala 282:24]
  reg [31:0] DMemory_394; // @[cpu.scala 282:24]
  reg [31:0] DMemory_395; // @[cpu.scala 282:24]
  reg [31:0] DMemory_396; // @[cpu.scala 282:24]
  reg [31:0] DMemory_397; // @[cpu.scala 282:24]
  reg [31:0] DMemory_398; // @[cpu.scala 282:24]
  reg [31:0] DMemory_399; // @[cpu.scala 282:24]
  reg [31:0] DMemory_400; // @[cpu.scala 282:24]
  reg [31:0] DMemory_401; // @[cpu.scala 282:24]
  reg [31:0] DMemory_402; // @[cpu.scala 282:24]
  reg [31:0] DMemory_403; // @[cpu.scala 282:24]
  reg [31:0] DMemory_404; // @[cpu.scala 282:24]
  reg [31:0] DMemory_405; // @[cpu.scala 282:24]
  reg [31:0] DMemory_406; // @[cpu.scala 282:24]
  reg [31:0] DMemory_407; // @[cpu.scala 282:24]
  reg [31:0] DMemory_408; // @[cpu.scala 282:24]
  reg [31:0] DMemory_409; // @[cpu.scala 282:24]
  reg [31:0] DMemory_410; // @[cpu.scala 282:24]
  reg [31:0] DMemory_411; // @[cpu.scala 282:24]
  reg [31:0] DMemory_412; // @[cpu.scala 282:24]
  reg [31:0] DMemory_413; // @[cpu.scala 282:24]
  reg [31:0] DMemory_414; // @[cpu.scala 282:24]
  reg [31:0] DMemory_415; // @[cpu.scala 282:24]
  reg [31:0] DMemory_416; // @[cpu.scala 282:24]
  reg [31:0] DMemory_417; // @[cpu.scala 282:24]
  reg [31:0] DMemory_418; // @[cpu.scala 282:24]
  reg [31:0] DMemory_419; // @[cpu.scala 282:24]
  reg [31:0] DMemory_420; // @[cpu.scala 282:24]
  reg [31:0] DMemory_421; // @[cpu.scala 282:24]
  reg [31:0] DMemory_422; // @[cpu.scala 282:24]
  reg [31:0] DMemory_423; // @[cpu.scala 282:24]
  reg [31:0] DMemory_424; // @[cpu.scala 282:24]
  reg [31:0] DMemory_425; // @[cpu.scala 282:24]
  reg [31:0] DMemory_426; // @[cpu.scala 282:24]
  reg [31:0] DMemory_427; // @[cpu.scala 282:24]
  reg [31:0] DMemory_428; // @[cpu.scala 282:24]
  reg [31:0] DMemory_429; // @[cpu.scala 282:24]
  reg [31:0] DMemory_430; // @[cpu.scala 282:24]
  reg [31:0] DMemory_431; // @[cpu.scala 282:24]
  reg [31:0] DMemory_432; // @[cpu.scala 282:24]
  reg [31:0] DMemory_433; // @[cpu.scala 282:24]
  reg [31:0] DMemory_434; // @[cpu.scala 282:24]
  reg [31:0] DMemory_435; // @[cpu.scala 282:24]
  reg [31:0] DMemory_436; // @[cpu.scala 282:24]
  reg [31:0] DMemory_437; // @[cpu.scala 282:24]
  reg [31:0] DMemory_438; // @[cpu.scala 282:24]
  reg [31:0] DMemory_439; // @[cpu.scala 282:24]
  reg [31:0] DMemory_440; // @[cpu.scala 282:24]
  reg [31:0] DMemory_441; // @[cpu.scala 282:24]
  reg [31:0] DMemory_442; // @[cpu.scala 282:24]
  reg [31:0] DMemory_443; // @[cpu.scala 282:24]
  reg [31:0] DMemory_444; // @[cpu.scala 282:24]
  reg [31:0] DMemory_445; // @[cpu.scala 282:24]
  reg [31:0] DMemory_446; // @[cpu.scala 282:24]
  reg [31:0] DMemory_447; // @[cpu.scala 282:24]
  reg [31:0] DMemory_448; // @[cpu.scala 282:24]
  reg [31:0] DMemory_449; // @[cpu.scala 282:24]
  reg [31:0] DMemory_450; // @[cpu.scala 282:24]
  reg [31:0] DMemory_451; // @[cpu.scala 282:24]
  reg [31:0] DMemory_452; // @[cpu.scala 282:24]
  reg [31:0] DMemory_453; // @[cpu.scala 282:24]
  reg [31:0] DMemory_454; // @[cpu.scala 282:24]
  reg [31:0] DMemory_455; // @[cpu.scala 282:24]
  reg [31:0] DMemory_456; // @[cpu.scala 282:24]
  reg [31:0] DMemory_457; // @[cpu.scala 282:24]
  reg [31:0] DMemory_458; // @[cpu.scala 282:24]
  reg [31:0] DMemory_459; // @[cpu.scala 282:24]
  reg [31:0] DMemory_460; // @[cpu.scala 282:24]
  reg [31:0] DMemory_461; // @[cpu.scala 282:24]
  reg [31:0] DMemory_462; // @[cpu.scala 282:24]
  reg [31:0] DMemory_463; // @[cpu.scala 282:24]
  reg [31:0] DMemory_464; // @[cpu.scala 282:24]
  reg [31:0] DMemory_465; // @[cpu.scala 282:24]
  reg [31:0] DMemory_466; // @[cpu.scala 282:24]
  reg [31:0] DMemory_467; // @[cpu.scala 282:24]
  reg [31:0] DMemory_468; // @[cpu.scala 282:24]
  reg [31:0] DMemory_469; // @[cpu.scala 282:24]
  reg [31:0] DMemory_470; // @[cpu.scala 282:24]
  reg [31:0] DMemory_471; // @[cpu.scala 282:24]
  reg [31:0] DMemory_472; // @[cpu.scala 282:24]
  reg [31:0] DMemory_473; // @[cpu.scala 282:24]
  reg [31:0] DMemory_474; // @[cpu.scala 282:24]
  reg [31:0] DMemory_475; // @[cpu.scala 282:24]
  reg [31:0] DMemory_476; // @[cpu.scala 282:24]
  reg [31:0] DMemory_477; // @[cpu.scala 282:24]
  reg [31:0] DMemory_478; // @[cpu.scala 282:24]
  reg [31:0] DMemory_479; // @[cpu.scala 282:24]
  reg [31:0] DMemory_480; // @[cpu.scala 282:24]
  reg [31:0] DMemory_481; // @[cpu.scala 282:24]
  reg [31:0] DMemory_482; // @[cpu.scala 282:24]
  reg [31:0] DMemory_483; // @[cpu.scala 282:24]
  reg [31:0] DMemory_484; // @[cpu.scala 282:24]
  reg [31:0] DMemory_485; // @[cpu.scala 282:24]
  reg [31:0] DMemory_486; // @[cpu.scala 282:24]
  reg [31:0] DMemory_487; // @[cpu.scala 282:24]
  reg [31:0] DMemory_488; // @[cpu.scala 282:24]
  reg [31:0] DMemory_489; // @[cpu.scala 282:24]
  reg [31:0] DMemory_490; // @[cpu.scala 282:24]
  reg [31:0] DMemory_491; // @[cpu.scala 282:24]
  reg [31:0] DMemory_492; // @[cpu.scala 282:24]
  reg [31:0] DMemory_493; // @[cpu.scala 282:24]
  reg [31:0] DMemory_494; // @[cpu.scala 282:24]
  reg [31:0] DMemory_495; // @[cpu.scala 282:24]
  reg [31:0] DMemory_496; // @[cpu.scala 282:24]
  reg [31:0] DMemory_497; // @[cpu.scala 282:24]
  reg [31:0] DMemory_498; // @[cpu.scala 282:24]
  reg [31:0] DMemory_499; // @[cpu.scala 282:24]
  reg [31:0] DMemory_500; // @[cpu.scala 282:24]
  reg [31:0] DMemory_501; // @[cpu.scala 282:24]
  reg [31:0] DMemory_502; // @[cpu.scala 282:24]
  reg [31:0] DMemory_503; // @[cpu.scala 282:24]
  reg [31:0] DMemory_504; // @[cpu.scala 282:24]
  reg [31:0] DMemory_505; // @[cpu.scala 282:24]
  reg [31:0] DMemory_506; // @[cpu.scala 282:24]
  reg [31:0] DMemory_507; // @[cpu.scala 282:24]
  reg [31:0] DMemory_508; // @[cpu.scala 282:24]
  reg [31:0] DMemory_509; // @[cpu.scala 282:24]
  reg [31:0] DMemory_510; // @[cpu.scala 282:24]
  reg [31:0] DMemory_511; // @[cpu.scala 282:24]
  reg [31:0] DMemory_512; // @[cpu.scala 282:24]
  reg [31:0] DMemory_513; // @[cpu.scala 282:24]
  reg [31:0] DMemory_514; // @[cpu.scala 282:24]
  reg [31:0] DMemory_515; // @[cpu.scala 282:24]
  reg [31:0] DMemory_516; // @[cpu.scala 282:24]
  reg [31:0] DMemory_517; // @[cpu.scala 282:24]
  reg [31:0] DMemory_518; // @[cpu.scala 282:24]
  reg [31:0] DMemory_519; // @[cpu.scala 282:24]
  reg [31:0] DMemory_520; // @[cpu.scala 282:24]
  reg [31:0] DMemory_521; // @[cpu.scala 282:24]
  reg [31:0] DMemory_522; // @[cpu.scala 282:24]
  reg [31:0] DMemory_523; // @[cpu.scala 282:24]
  reg [31:0] DMemory_524; // @[cpu.scala 282:24]
  reg [31:0] DMemory_525; // @[cpu.scala 282:24]
  reg [31:0] DMemory_526; // @[cpu.scala 282:24]
  reg [31:0] DMemory_527; // @[cpu.scala 282:24]
  reg [31:0] DMemory_528; // @[cpu.scala 282:24]
  reg [31:0] DMemory_529; // @[cpu.scala 282:24]
  reg [31:0] DMemory_530; // @[cpu.scala 282:24]
  reg [31:0] DMemory_531; // @[cpu.scala 282:24]
  reg [31:0] DMemory_532; // @[cpu.scala 282:24]
  reg [31:0] DMemory_533; // @[cpu.scala 282:24]
  reg [31:0] DMemory_534; // @[cpu.scala 282:24]
  reg [31:0] DMemory_535; // @[cpu.scala 282:24]
  reg [31:0] DMemory_536; // @[cpu.scala 282:24]
  reg [31:0] DMemory_537; // @[cpu.scala 282:24]
  reg [31:0] DMemory_538; // @[cpu.scala 282:24]
  reg [31:0] DMemory_539; // @[cpu.scala 282:24]
  reg [31:0] DMemory_540; // @[cpu.scala 282:24]
  reg [31:0] DMemory_541; // @[cpu.scala 282:24]
  reg [31:0] DMemory_542; // @[cpu.scala 282:24]
  reg [31:0] DMemory_543; // @[cpu.scala 282:24]
  reg [31:0] DMemory_544; // @[cpu.scala 282:24]
  reg [31:0] DMemory_545; // @[cpu.scala 282:24]
  reg [31:0] DMemory_546; // @[cpu.scala 282:24]
  reg [31:0] DMemory_547; // @[cpu.scala 282:24]
  reg [31:0] DMemory_548; // @[cpu.scala 282:24]
  reg [31:0] DMemory_549; // @[cpu.scala 282:24]
  reg [31:0] DMemory_550; // @[cpu.scala 282:24]
  reg [31:0] DMemory_551; // @[cpu.scala 282:24]
  reg [31:0] DMemory_552; // @[cpu.scala 282:24]
  reg [31:0] DMemory_553; // @[cpu.scala 282:24]
  reg [31:0] DMemory_554; // @[cpu.scala 282:24]
  reg [31:0] DMemory_555; // @[cpu.scala 282:24]
  reg [31:0] DMemory_556; // @[cpu.scala 282:24]
  reg [31:0] DMemory_557; // @[cpu.scala 282:24]
  reg [31:0] DMemory_558; // @[cpu.scala 282:24]
  reg [31:0] DMemory_559; // @[cpu.scala 282:24]
  reg [31:0] DMemory_560; // @[cpu.scala 282:24]
  reg [31:0] DMemory_561; // @[cpu.scala 282:24]
  reg [31:0] DMemory_562; // @[cpu.scala 282:24]
  reg [31:0] DMemory_563; // @[cpu.scala 282:24]
  reg [31:0] DMemory_564; // @[cpu.scala 282:24]
  reg [31:0] DMemory_565; // @[cpu.scala 282:24]
  reg [31:0] DMemory_566; // @[cpu.scala 282:24]
  reg [31:0] DMemory_567; // @[cpu.scala 282:24]
  reg [31:0] DMemory_568; // @[cpu.scala 282:24]
  reg [31:0] DMemory_569; // @[cpu.scala 282:24]
  reg [31:0] DMemory_570; // @[cpu.scala 282:24]
  reg [31:0] DMemory_571; // @[cpu.scala 282:24]
  reg [31:0] DMemory_572; // @[cpu.scala 282:24]
  reg [31:0] DMemory_573; // @[cpu.scala 282:24]
  reg [31:0] DMemory_574; // @[cpu.scala 282:24]
  reg [31:0] DMemory_575; // @[cpu.scala 282:24]
  reg [31:0] DMemory_576; // @[cpu.scala 282:24]
  reg [31:0] DMemory_577; // @[cpu.scala 282:24]
  reg [31:0] DMemory_578; // @[cpu.scala 282:24]
  reg [31:0] DMemory_579; // @[cpu.scala 282:24]
  reg [31:0] DMemory_580; // @[cpu.scala 282:24]
  reg [31:0] DMemory_581; // @[cpu.scala 282:24]
  reg [31:0] DMemory_582; // @[cpu.scala 282:24]
  reg [31:0] DMemory_583; // @[cpu.scala 282:24]
  reg [31:0] DMemory_584; // @[cpu.scala 282:24]
  reg [31:0] DMemory_585; // @[cpu.scala 282:24]
  reg [31:0] DMemory_586; // @[cpu.scala 282:24]
  reg [31:0] DMemory_587; // @[cpu.scala 282:24]
  reg [31:0] DMemory_588; // @[cpu.scala 282:24]
  reg [31:0] DMemory_589; // @[cpu.scala 282:24]
  reg [31:0] DMemory_590; // @[cpu.scala 282:24]
  reg [31:0] DMemory_591; // @[cpu.scala 282:24]
  reg [31:0] DMemory_592; // @[cpu.scala 282:24]
  reg [31:0] DMemory_593; // @[cpu.scala 282:24]
  reg [31:0] DMemory_594; // @[cpu.scala 282:24]
  reg [31:0] DMemory_595; // @[cpu.scala 282:24]
  reg [31:0] DMemory_596; // @[cpu.scala 282:24]
  reg [31:0] DMemory_597; // @[cpu.scala 282:24]
  reg [31:0] DMemory_598; // @[cpu.scala 282:24]
  reg [31:0] DMemory_599; // @[cpu.scala 282:24]
  reg [31:0] DMemory_600; // @[cpu.scala 282:24]
  reg [31:0] DMemory_601; // @[cpu.scala 282:24]
  reg [31:0] DMemory_602; // @[cpu.scala 282:24]
  reg [31:0] DMemory_603; // @[cpu.scala 282:24]
  reg [31:0] DMemory_604; // @[cpu.scala 282:24]
  reg [31:0] DMemory_605; // @[cpu.scala 282:24]
  reg [31:0] DMemory_606; // @[cpu.scala 282:24]
  reg [31:0] DMemory_607; // @[cpu.scala 282:24]
  reg [31:0] DMemory_608; // @[cpu.scala 282:24]
  reg [31:0] DMemory_609; // @[cpu.scala 282:24]
  reg [31:0] DMemory_610; // @[cpu.scala 282:24]
  reg [31:0] DMemory_611; // @[cpu.scala 282:24]
  reg [31:0] DMemory_612; // @[cpu.scala 282:24]
  reg [31:0] DMemory_613; // @[cpu.scala 282:24]
  reg [31:0] DMemory_614; // @[cpu.scala 282:24]
  reg [31:0] DMemory_615; // @[cpu.scala 282:24]
  reg [31:0] DMemory_616; // @[cpu.scala 282:24]
  reg [31:0] DMemory_617; // @[cpu.scala 282:24]
  reg [31:0] DMemory_618; // @[cpu.scala 282:24]
  reg [31:0] DMemory_619; // @[cpu.scala 282:24]
  reg [31:0] DMemory_620; // @[cpu.scala 282:24]
  reg [31:0] DMemory_621; // @[cpu.scala 282:24]
  reg [31:0] DMemory_622; // @[cpu.scala 282:24]
  reg [31:0] DMemory_623; // @[cpu.scala 282:24]
  reg [31:0] DMemory_624; // @[cpu.scala 282:24]
  reg [31:0] DMemory_625; // @[cpu.scala 282:24]
  reg [31:0] DMemory_626; // @[cpu.scala 282:24]
  reg [31:0] DMemory_627; // @[cpu.scala 282:24]
  reg [31:0] DMemory_628; // @[cpu.scala 282:24]
  reg [31:0] DMemory_629; // @[cpu.scala 282:24]
  reg [31:0] DMemory_630; // @[cpu.scala 282:24]
  reg [31:0] DMemory_631; // @[cpu.scala 282:24]
  reg [31:0] DMemory_632; // @[cpu.scala 282:24]
  reg [31:0] DMemory_633; // @[cpu.scala 282:24]
  reg [31:0] DMemory_634; // @[cpu.scala 282:24]
  reg [31:0] DMemory_635; // @[cpu.scala 282:24]
  reg [31:0] DMemory_636; // @[cpu.scala 282:24]
  reg [31:0] DMemory_637; // @[cpu.scala 282:24]
  reg [31:0] DMemory_638; // @[cpu.scala 282:24]
  reg [31:0] DMemory_639; // @[cpu.scala 282:24]
  reg [31:0] DMemory_640; // @[cpu.scala 282:24]
  reg [31:0] DMemory_641; // @[cpu.scala 282:24]
  reg [31:0] DMemory_642; // @[cpu.scala 282:24]
  reg [31:0] DMemory_643; // @[cpu.scala 282:24]
  reg [31:0] DMemory_644; // @[cpu.scala 282:24]
  reg [31:0] DMemory_645; // @[cpu.scala 282:24]
  reg [31:0] DMemory_646; // @[cpu.scala 282:24]
  reg [31:0] DMemory_647; // @[cpu.scala 282:24]
  reg [31:0] DMemory_648; // @[cpu.scala 282:24]
  reg [31:0] DMemory_649; // @[cpu.scala 282:24]
  reg [31:0] DMemory_650; // @[cpu.scala 282:24]
  reg [31:0] DMemory_651; // @[cpu.scala 282:24]
  reg [31:0] DMemory_652; // @[cpu.scala 282:24]
  reg [31:0] DMemory_653; // @[cpu.scala 282:24]
  reg [31:0] DMemory_654; // @[cpu.scala 282:24]
  reg [31:0] DMemory_655; // @[cpu.scala 282:24]
  reg [31:0] DMemory_656; // @[cpu.scala 282:24]
  reg [31:0] DMemory_657; // @[cpu.scala 282:24]
  reg [31:0] DMemory_658; // @[cpu.scala 282:24]
  reg [31:0] DMemory_659; // @[cpu.scala 282:24]
  reg [31:0] DMemory_660; // @[cpu.scala 282:24]
  reg [31:0] DMemory_661; // @[cpu.scala 282:24]
  reg [31:0] DMemory_662; // @[cpu.scala 282:24]
  reg [31:0] DMemory_663; // @[cpu.scala 282:24]
  reg [31:0] DMemory_664; // @[cpu.scala 282:24]
  reg [31:0] DMemory_665; // @[cpu.scala 282:24]
  reg [31:0] DMemory_666; // @[cpu.scala 282:24]
  reg [31:0] DMemory_667; // @[cpu.scala 282:24]
  reg [31:0] DMemory_668; // @[cpu.scala 282:24]
  reg [31:0] DMemory_669; // @[cpu.scala 282:24]
  reg [31:0] DMemory_670; // @[cpu.scala 282:24]
  reg [31:0] DMemory_671; // @[cpu.scala 282:24]
  reg [31:0] DMemory_672; // @[cpu.scala 282:24]
  reg [31:0] DMemory_673; // @[cpu.scala 282:24]
  reg [31:0] DMemory_674; // @[cpu.scala 282:24]
  reg [31:0] DMemory_675; // @[cpu.scala 282:24]
  reg [31:0] DMemory_676; // @[cpu.scala 282:24]
  reg [31:0] DMemory_677; // @[cpu.scala 282:24]
  reg [31:0] DMemory_678; // @[cpu.scala 282:24]
  reg [31:0] DMemory_679; // @[cpu.scala 282:24]
  reg [31:0] DMemory_680; // @[cpu.scala 282:24]
  reg [31:0] DMemory_681; // @[cpu.scala 282:24]
  reg [31:0] DMemory_682; // @[cpu.scala 282:24]
  reg [31:0] DMemory_683; // @[cpu.scala 282:24]
  reg [31:0] DMemory_684; // @[cpu.scala 282:24]
  reg [31:0] DMemory_685; // @[cpu.scala 282:24]
  reg [31:0] DMemory_686; // @[cpu.scala 282:24]
  reg [31:0] DMemory_687; // @[cpu.scala 282:24]
  reg [31:0] DMemory_688; // @[cpu.scala 282:24]
  reg [31:0] DMemory_689; // @[cpu.scala 282:24]
  reg [31:0] DMemory_690; // @[cpu.scala 282:24]
  reg [31:0] DMemory_691; // @[cpu.scala 282:24]
  reg [31:0] DMemory_692; // @[cpu.scala 282:24]
  reg [31:0] DMemory_693; // @[cpu.scala 282:24]
  reg [31:0] DMemory_694; // @[cpu.scala 282:24]
  reg [31:0] DMemory_695; // @[cpu.scala 282:24]
  reg [31:0] DMemory_696; // @[cpu.scala 282:24]
  reg [31:0] DMemory_697; // @[cpu.scala 282:24]
  reg [31:0] DMemory_698; // @[cpu.scala 282:24]
  reg [31:0] DMemory_699; // @[cpu.scala 282:24]
  reg [31:0] DMemory_700; // @[cpu.scala 282:24]
  reg [31:0] DMemory_701; // @[cpu.scala 282:24]
  reg [31:0] DMemory_702; // @[cpu.scala 282:24]
  reg [31:0] DMemory_703; // @[cpu.scala 282:24]
  reg [31:0] DMemory_704; // @[cpu.scala 282:24]
  reg [31:0] DMemory_705; // @[cpu.scala 282:24]
  reg [31:0] DMemory_706; // @[cpu.scala 282:24]
  reg [31:0] DMemory_707; // @[cpu.scala 282:24]
  reg [31:0] DMemory_708; // @[cpu.scala 282:24]
  reg [31:0] DMemory_709; // @[cpu.scala 282:24]
  reg [31:0] DMemory_710; // @[cpu.scala 282:24]
  reg [31:0] DMemory_711; // @[cpu.scala 282:24]
  reg [31:0] DMemory_712; // @[cpu.scala 282:24]
  reg [31:0] DMemory_713; // @[cpu.scala 282:24]
  reg [31:0] DMemory_714; // @[cpu.scala 282:24]
  reg [31:0] DMemory_715; // @[cpu.scala 282:24]
  reg [31:0] DMemory_716; // @[cpu.scala 282:24]
  reg [31:0] DMemory_717; // @[cpu.scala 282:24]
  reg [31:0] DMemory_718; // @[cpu.scala 282:24]
  reg [31:0] DMemory_719; // @[cpu.scala 282:24]
  reg [31:0] DMemory_720; // @[cpu.scala 282:24]
  reg [31:0] DMemory_721; // @[cpu.scala 282:24]
  reg [31:0] DMemory_722; // @[cpu.scala 282:24]
  reg [31:0] DMemory_723; // @[cpu.scala 282:24]
  reg [31:0] DMemory_724; // @[cpu.scala 282:24]
  reg [31:0] DMemory_725; // @[cpu.scala 282:24]
  reg [31:0] DMemory_726; // @[cpu.scala 282:24]
  reg [31:0] DMemory_727; // @[cpu.scala 282:24]
  reg [31:0] DMemory_728; // @[cpu.scala 282:24]
  reg [31:0] DMemory_729; // @[cpu.scala 282:24]
  reg [31:0] DMemory_730; // @[cpu.scala 282:24]
  reg [31:0] DMemory_731; // @[cpu.scala 282:24]
  reg [31:0] DMemory_732; // @[cpu.scala 282:24]
  reg [31:0] DMemory_733; // @[cpu.scala 282:24]
  reg [31:0] DMemory_734; // @[cpu.scala 282:24]
  reg [31:0] DMemory_735; // @[cpu.scala 282:24]
  reg [31:0] DMemory_736; // @[cpu.scala 282:24]
  reg [31:0] DMemory_737; // @[cpu.scala 282:24]
  reg [31:0] DMemory_738; // @[cpu.scala 282:24]
  reg [31:0] DMemory_739; // @[cpu.scala 282:24]
  reg [31:0] DMemory_740; // @[cpu.scala 282:24]
  reg [31:0] DMemory_741; // @[cpu.scala 282:24]
  reg [31:0] DMemory_742; // @[cpu.scala 282:24]
  reg [31:0] DMemory_743; // @[cpu.scala 282:24]
  reg [31:0] DMemory_744; // @[cpu.scala 282:24]
  reg [31:0] DMemory_745; // @[cpu.scala 282:24]
  reg [31:0] DMemory_746; // @[cpu.scala 282:24]
  reg [31:0] DMemory_747; // @[cpu.scala 282:24]
  reg [31:0] DMemory_748; // @[cpu.scala 282:24]
  reg [31:0] DMemory_749; // @[cpu.scala 282:24]
  reg [31:0] DMemory_750; // @[cpu.scala 282:24]
  reg [31:0] DMemory_751; // @[cpu.scala 282:24]
  reg [31:0] DMemory_752; // @[cpu.scala 282:24]
  reg [31:0] DMemory_753; // @[cpu.scala 282:24]
  reg [31:0] DMemory_754; // @[cpu.scala 282:24]
  reg [31:0] DMemory_755; // @[cpu.scala 282:24]
  reg [31:0] DMemory_756; // @[cpu.scala 282:24]
  reg [31:0] DMemory_757; // @[cpu.scala 282:24]
  reg [31:0] DMemory_758; // @[cpu.scala 282:24]
  reg [31:0] DMemory_759; // @[cpu.scala 282:24]
  reg [31:0] DMemory_760; // @[cpu.scala 282:24]
  reg [31:0] DMemory_761; // @[cpu.scala 282:24]
  reg [31:0] DMemory_762; // @[cpu.scala 282:24]
  reg [31:0] DMemory_763; // @[cpu.scala 282:24]
  reg [31:0] DMemory_764; // @[cpu.scala 282:24]
  reg [31:0] DMemory_765; // @[cpu.scala 282:24]
  reg [31:0] DMemory_766; // @[cpu.scala 282:24]
  reg [31:0] DMemory_767; // @[cpu.scala 282:24]
  reg [31:0] DMemory_768; // @[cpu.scala 282:24]
  reg [31:0] DMemory_769; // @[cpu.scala 282:24]
  reg [31:0] DMemory_770; // @[cpu.scala 282:24]
  reg [31:0] DMemory_771; // @[cpu.scala 282:24]
  reg [31:0] DMemory_772; // @[cpu.scala 282:24]
  reg [31:0] DMemory_773; // @[cpu.scala 282:24]
  reg [31:0] DMemory_774; // @[cpu.scala 282:24]
  reg [31:0] DMemory_775; // @[cpu.scala 282:24]
  reg [31:0] DMemory_776; // @[cpu.scala 282:24]
  reg [31:0] DMemory_777; // @[cpu.scala 282:24]
  reg [31:0] DMemory_778; // @[cpu.scala 282:24]
  reg [31:0] DMemory_779; // @[cpu.scala 282:24]
  reg [31:0] DMemory_780; // @[cpu.scala 282:24]
  reg [31:0] DMemory_781; // @[cpu.scala 282:24]
  reg [31:0] DMemory_782; // @[cpu.scala 282:24]
  reg [31:0] DMemory_783; // @[cpu.scala 282:24]
  reg [31:0] DMemory_784; // @[cpu.scala 282:24]
  reg [31:0] DMemory_785; // @[cpu.scala 282:24]
  reg [31:0] DMemory_786; // @[cpu.scala 282:24]
  reg [31:0] DMemory_787; // @[cpu.scala 282:24]
  reg [31:0] DMemory_788; // @[cpu.scala 282:24]
  reg [31:0] DMemory_789; // @[cpu.scala 282:24]
  reg [31:0] DMemory_790; // @[cpu.scala 282:24]
  reg [31:0] DMemory_791; // @[cpu.scala 282:24]
  reg [31:0] DMemory_792; // @[cpu.scala 282:24]
  reg [31:0] DMemory_793; // @[cpu.scala 282:24]
  reg [31:0] DMemory_794; // @[cpu.scala 282:24]
  reg [31:0] DMemory_795; // @[cpu.scala 282:24]
  reg [31:0] DMemory_796; // @[cpu.scala 282:24]
  reg [31:0] DMemory_797; // @[cpu.scala 282:24]
  reg [31:0] DMemory_798; // @[cpu.scala 282:24]
  reg [31:0] DMemory_799; // @[cpu.scala 282:24]
  reg [31:0] DMemory_800; // @[cpu.scala 282:24]
  reg [31:0] DMemory_801; // @[cpu.scala 282:24]
  reg [31:0] DMemory_802; // @[cpu.scala 282:24]
  reg [31:0] DMemory_803; // @[cpu.scala 282:24]
  reg [31:0] DMemory_804; // @[cpu.scala 282:24]
  reg [31:0] DMemory_805; // @[cpu.scala 282:24]
  reg [31:0] DMemory_806; // @[cpu.scala 282:24]
  reg [31:0] DMemory_807; // @[cpu.scala 282:24]
  reg [31:0] DMemory_808; // @[cpu.scala 282:24]
  reg [31:0] DMemory_809; // @[cpu.scala 282:24]
  reg [31:0] DMemory_810; // @[cpu.scala 282:24]
  reg [31:0] DMemory_811; // @[cpu.scala 282:24]
  reg [31:0] DMemory_812; // @[cpu.scala 282:24]
  reg [31:0] DMemory_813; // @[cpu.scala 282:24]
  reg [31:0] DMemory_814; // @[cpu.scala 282:24]
  reg [31:0] DMemory_815; // @[cpu.scala 282:24]
  reg [31:0] DMemory_816; // @[cpu.scala 282:24]
  reg [31:0] DMemory_817; // @[cpu.scala 282:24]
  reg [31:0] DMemory_818; // @[cpu.scala 282:24]
  reg [31:0] DMemory_819; // @[cpu.scala 282:24]
  reg [31:0] DMemory_820; // @[cpu.scala 282:24]
  reg [31:0] DMemory_821; // @[cpu.scala 282:24]
  reg [31:0] DMemory_822; // @[cpu.scala 282:24]
  reg [31:0] DMemory_823; // @[cpu.scala 282:24]
  reg [31:0] DMemory_824; // @[cpu.scala 282:24]
  reg [31:0] DMemory_825; // @[cpu.scala 282:24]
  reg [31:0] DMemory_826; // @[cpu.scala 282:24]
  reg [31:0] DMemory_827; // @[cpu.scala 282:24]
  reg [31:0] DMemory_828; // @[cpu.scala 282:24]
  reg [31:0] DMemory_829; // @[cpu.scala 282:24]
  reg [31:0] DMemory_830; // @[cpu.scala 282:24]
  reg [31:0] DMemory_831; // @[cpu.scala 282:24]
  reg [31:0] DMemory_832; // @[cpu.scala 282:24]
  reg [31:0] DMemory_833; // @[cpu.scala 282:24]
  reg [31:0] DMemory_834; // @[cpu.scala 282:24]
  reg [31:0] DMemory_835; // @[cpu.scala 282:24]
  reg [31:0] DMemory_836; // @[cpu.scala 282:24]
  reg [31:0] DMemory_837; // @[cpu.scala 282:24]
  reg [31:0] DMemory_838; // @[cpu.scala 282:24]
  reg [31:0] DMemory_839; // @[cpu.scala 282:24]
  reg [31:0] DMemory_840; // @[cpu.scala 282:24]
  reg [31:0] DMemory_841; // @[cpu.scala 282:24]
  reg [31:0] DMemory_842; // @[cpu.scala 282:24]
  reg [31:0] DMemory_843; // @[cpu.scala 282:24]
  reg [31:0] DMemory_844; // @[cpu.scala 282:24]
  reg [31:0] DMemory_845; // @[cpu.scala 282:24]
  reg [31:0] DMemory_846; // @[cpu.scala 282:24]
  reg [31:0] DMemory_847; // @[cpu.scala 282:24]
  reg [31:0] DMemory_848; // @[cpu.scala 282:24]
  reg [31:0] DMemory_849; // @[cpu.scala 282:24]
  reg [31:0] DMemory_850; // @[cpu.scala 282:24]
  reg [31:0] DMemory_851; // @[cpu.scala 282:24]
  reg [31:0] DMemory_852; // @[cpu.scala 282:24]
  reg [31:0] DMemory_853; // @[cpu.scala 282:24]
  reg [31:0] DMemory_854; // @[cpu.scala 282:24]
  reg [31:0] DMemory_855; // @[cpu.scala 282:24]
  reg [31:0] DMemory_856; // @[cpu.scala 282:24]
  reg [31:0] DMemory_857; // @[cpu.scala 282:24]
  reg [31:0] DMemory_858; // @[cpu.scala 282:24]
  reg [31:0] DMemory_859; // @[cpu.scala 282:24]
  reg [31:0] DMemory_860; // @[cpu.scala 282:24]
  reg [31:0] DMemory_861; // @[cpu.scala 282:24]
  reg [31:0] DMemory_862; // @[cpu.scala 282:24]
  reg [31:0] DMemory_863; // @[cpu.scala 282:24]
  reg [31:0] DMemory_864; // @[cpu.scala 282:24]
  reg [31:0] DMemory_865; // @[cpu.scala 282:24]
  reg [31:0] DMemory_866; // @[cpu.scala 282:24]
  reg [31:0] DMemory_867; // @[cpu.scala 282:24]
  reg [31:0] DMemory_868; // @[cpu.scala 282:24]
  reg [31:0] DMemory_869; // @[cpu.scala 282:24]
  reg [31:0] DMemory_870; // @[cpu.scala 282:24]
  reg [31:0] DMemory_871; // @[cpu.scala 282:24]
  reg [31:0] DMemory_872; // @[cpu.scala 282:24]
  reg [31:0] DMemory_873; // @[cpu.scala 282:24]
  reg [31:0] DMemory_874; // @[cpu.scala 282:24]
  reg [31:0] DMemory_875; // @[cpu.scala 282:24]
  reg [31:0] DMemory_876; // @[cpu.scala 282:24]
  reg [31:0] DMemory_877; // @[cpu.scala 282:24]
  reg [31:0] DMemory_878; // @[cpu.scala 282:24]
  reg [31:0] DMemory_879; // @[cpu.scala 282:24]
  reg [31:0] DMemory_880; // @[cpu.scala 282:24]
  reg [31:0] DMemory_881; // @[cpu.scala 282:24]
  reg [31:0] DMemory_882; // @[cpu.scala 282:24]
  reg [31:0] DMemory_883; // @[cpu.scala 282:24]
  reg [31:0] DMemory_884; // @[cpu.scala 282:24]
  reg [31:0] DMemory_885; // @[cpu.scala 282:24]
  reg [31:0] DMemory_886; // @[cpu.scala 282:24]
  reg [31:0] DMemory_887; // @[cpu.scala 282:24]
  reg [31:0] DMemory_888; // @[cpu.scala 282:24]
  reg [31:0] DMemory_889; // @[cpu.scala 282:24]
  reg [31:0] DMemory_890; // @[cpu.scala 282:24]
  reg [31:0] DMemory_891; // @[cpu.scala 282:24]
  reg [31:0] DMemory_892; // @[cpu.scala 282:24]
  reg [31:0] DMemory_893; // @[cpu.scala 282:24]
  reg [31:0] DMemory_894; // @[cpu.scala 282:24]
  reg [31:0] DMemory_895; // @[cpu.scala 282:24]
  reg [31:0] DMemory_896; // @[cpu.scala 282:24]
  reg [31:0] DMemory_897; // @[cpu.scala 282:24]
  reg [31:0] DMemory_898; // @[cpu.scala 282:24]
  reg [31:0] DMemory_899; // @[cpu.scala 282:24]
  reg [31:0] DMemory_900; // @[cpu.scala 282:24]
  reg [31:0] DMemory_901; // @[cpu.scala 282:24]
  reg [31:0] DMemory_902; // @[cpu.scala 282:24]
  reg [31:0] DMemory_903; // @[cpu.scala 282:24]
  reg [31:0] DMemory_904; // @[cpu.scala 282:24]
  reg [31:0] DMemory_905; // @[cpu.scala 282:24]
  reg [31:0] DMemory_906; // @[cpu.scala 282:24]
  reg [31:0] DMemory_907; // @[cpu.scala 282:24]
  reg [31:0] DMemory_908; // @[cpu.scala 282:24]
  reg [31:0] DMemory_909; // @[cpu.scala 282:24]
  reg [31:0] DMemory_910; // @[cpu.scala 282:24]
  reg [31:0] DMemory_911; // @[cpu.scala 282:24]
  reg [31:0] DMemory_912; // @[cpu.scala 282:24]
  reg [31:0] DMemory_913; // @[cpu.scala 282:24]
  reg [31:0] DMemory_914; // @[cpu.scala 282:24]
  reg [31:0] DMemory_915; // @[cpu.scala 282:24]
  reg [31:0] DMemory_916; // @[cpu.scala 282:24]
  reg [31:0] DMemory_917; // @[cpu.scala 282:24]
  reg [31:0] DMemory_918; // @[cpu.scala 282:24]
  reg [31:0] DMemory_919; // @[cpu.scala 282:24]
  reg [31:0] DMemory_920; // @[cpu.scala 282:24]
  reg [31:0] DMemory_921; // @[cpu.scala 282:24]
  reg [31:0] DMemory_922; // @[cpu.scala 282:24]
  reg [31:0] DMemory_923; // @[cpu.scala 282:24]
  reg [31:0] DMemory_924; // @[cpu.scala 282:24]
  reg [31:0] DMemory_925; // @[cpu.scala 282:24]
  reg [31:0] DMemory_926; // @[cpu.scala 282:24]
  reg [31:0] DMemory_927; // @[cpu.scala 282:24]
  reg [31:0] DMemory_928; // @[cpu.scala 282:24]
  reg [31:0] DMemory_929; // @[cpu.scala 282:24]
  reg [31:0] DMemory_930; // @[cpu.scala 282:24]
  reg [31:0] DMemory_931; // @[cpu.scala 282:24]
  reg [31:0] DMemory_932; // @[cpu.scala 282:24]
  reg [31:0] DMemory_933; // @[cpu.scala 282:24]
  reg [31:0] DMemory_934; // @[cpu.scala 282:24]
  reg [31:0] DMemory_935; // @[cpu.scala 282:24]
  reg [31:0] DMemory_936; // @[cpu.scala 282:24]
  reg [31:0] DMemory_937; // @[cpu.scala 282:24]
  reg [31:0] DMemory_938; // @[cpu.scala 282:24]
  reg [31:0] DMemory_939; // @[cpu.scala 282:24]
  reg [31:0] DMemory_940; // @[cpu.scala 282:24]
  reg [31:0] DMemory_941; // @[cpu.scala 282:24]
  reg [31:0] DMemory_942; // @[cpu.scala 282:24]
  reg [31:0] DMemory_943; // @[cpu.scala 282:24]
  reg [31:0] DMemory_944; // @[cpu.scala 282:24]
  reg [31:0] DMemory_945; // @[cpu.scala 282:24]
  reg [31:0] DMemory_946; // @[cpu.scala 282:24]
  reg [31:0] DMemory_947; // @[cpu.scala 282:24]
  reg [31:0] DMemory_948; // @[cpu.scala 282:24]
  reg [31:0] DMemory_949; // @[cpu.scala 282:24]
  reg [31:0] DMemory_950; // @[cpu.scala 282:24]
  reg [31:0] DMemory_951; // @[cpu.scala 282:24]
  reg [31:0] DMemory_952; // @[cpu.scala 282:24]
  reg [31:0] DMemory_953; // @[cpu.scala 282:24]
  reg [31:0] DMemory_954; // @[cpu.scala 282:24]
  reg [31:0] DMemory_955; // @[cpu.scala 282:24]
  reg [31:0] DMemory_956; // @[cpu.scala 282:24]
  reg [31:0] DMemory_957; // @[cpu.scala 282:24]
  reg [31:0] DMemory_958; // @[cpu.scala 282:24]
  reg [31:0] DMemory_959; // @[cpu.scala 282:24]
  reg [31:0] DMemory_960; // @[cpu.scala 282:24]
  reg [31:0] DMemory_961; // @[cpu.scala 282:24]
  reg [31:0] DMemory_962; // @[cpu.scala 282:24]
  reg [31:0] DMemory_963; // @[cpu.scala 282:24]
  reg [31:0] DMemory_964; // @[cpu.scala 282:24]
  reg [31:0] DMemory_965; // @[cpu.scala 282:24]
  reg [31:0] DMemory_966; // @[cpu.scala 282:24]
  reg [31:0] DMemory_967; // @[cpu.scala 282:24]
  reg [31:0] DMemory_968; // @[cpu.scala 282:24]
  reg [31:0] DMemory_969; // @[cpu.scala 282:24]
  reg [31:0] DMemory_970; // @[cpu.scala 282:24]
  reg [31:0] DMemory_971; // @[cpu.scala 282:24]
  reg [31:0] DMemory_972; // @[cpu.scala 282:24]
  reg [31:0] DMemory_973; // @[cpu.scala 282:24]
  reg [31:0] DMemory_974; // @[cpu.scala 282:24]
  reg [31:0] DMemory_975; // @[cpu.scala 282:24]
  reg [31:0] DMemory_976; // @[cpu.scala 282:24]
  reg [31:0] DMemory_977; // @[cpu.scala 282:24]
  reg [31:0] DMemory_978; // @[cpu.scala 282:24]
  reg [31:0] DMemory_979; // @[cpu.scala 282:24]
  reg [31:0] DMemory_980; // @[cpu.scala 282:24]
  reg [31:0] DMemory_981; // @[cpu.scala 282:24]
  reg [31:0] DMemory_982; // @[cpu.scala 282:24]
  reg [31:0] DMemory_983; // @[cpu.scala 282:24]
  reg [31:0] DMemory_984; // @[cpu.scala 282:24]
  reg [31:0] DMemory_985; // @[cpu.scala 282:24]
  reg [31:0] DMemory_986; // @[cpu.scala 282:24]
  reg [31:0] DMemory_987; // @[cpu.scala 282:24]
  reg [31:0] DMemory_988; // @[cpu.scala 282:24]
  reg [31:0] DMemory_989; // @[cpu.scala 282:24]
  reg [31:0] DMemory_990; // @[cpu.scala 282:24]
  reg [31:0] DMemory_991; // @[cpu.scala 282:24]
  reg [31:0] DMemory_992; // @[cpu.scala 282:24]
  reg [31:0] DMemory_993; // @[cpu.scala 282:24]
  reg [31:0] DMemory_994; // @[cpu.scala 282:24]
  reg [31:0] DMemory_995; // @[cpu.scala 282:24]
  reg [31:0] DMemory_996; // @[cpu.scala 282:24]
  reg [31:0] DMemory_997; // @[cpu.scala 282:24]
  reg [31:0] DMemory_998; // @[cpu.scala 282:24]
  reg [31:0] DMemory_999; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1000; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1001; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1002; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1003; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1004; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1005; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1006; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1007; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1008; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1009; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1010; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1011; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1012; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1013; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1014; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1015; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1016; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1017; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1018; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1019; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1020; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1021; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1022; // @[cpu.scala 282:24]
  reg [31:0] DMemory_1023; // @[cpu.scala 282:24]
  reg [31:0] IMemory_0; // @[cpu.scala 283:24]
  reg [31:0] IMemory_1; // @[cpu.scala 283:24]
  reg [31:0] IFIDIR; // @[cpu.scala 286:49]
  reg [31:0] IDEXIR; // @[cpu.scala 286:49]
  reg [31:0] EXMEMIR; // @[cpu.scala 286:49]
  reg [31:0] MEMWBIR; // @[cpu.scala 286:49]
  reg [63:0] CurPC; // @[cpu.scala 289:22]
  wire [4:0] EXMEMrd = EXMEMIR[11:7]; // @[cpu.scala 321:32]
  wire [4:0] IDEXrd = IDEXIR[11:7]; // @[cpu.scala 322:30]
  wire [2:0] IFID_funct3 = IFIDIR[14:12]; // @[cpu.scala 323:29]
  wire [4:0] IFIDrs1 = io_rvfi_rst ? IFIDIR[19:15] : IFIDIR[19:15]; // @[cpu.scala 299:21 301:13 313:13]
  wire [4:0] MEMWBrd = io_rvfi_rst ? MEMWBIR[11:7] : MEMWBIR[11:7]; // @[cpu.scala 299:21 307:13 319:13]
  wire  _bypassAFromWB_T_1 = IFIDrs1 != 5'h0; // @[cpu.scala 326:41]
  wire [6:0] MEMWBop = io_rvfi_rst ? MEMWBIR[6:0] : MEMWBIR[6:0]; // @[cpu.scala 299:21 306:13 318:13]
  wire  _bypassAFromWB_T_3 = MEMWBop == 7'h33; // @[cpu.scala 326:62]
  wire  _bypassAFromWB_T_4 = MEMWBop == 7'h3; // @[cpu.scala 326:83]
  wire  _bypassAFromWB_T_5 = MEMWBop == 7'h33 | MEMWBop == 7'h3; // @[cpu.scala 326:72]
  wire  bypassAFromWB = IFIDrs1 == MEMWBrd & IFIDrs1 != 5'h0 & (MEMWBop == 7'h33 | MEMWBop == 7'h3); // @[cpu.scala 326:50]
  wire [4:0] IFIDrs2 = io_rvfi_rst ? IFIDIR[24:20] : IFIDIR[24:20]; // @[cpu.scala 299:21 302:13 314:13]
  wire  _bypassBFromWB_T_1 = IFIDrs2 != 5'h0; // @[cpu.scala 328:41]
  wire  bypassBFromWB = IFIDrs2 == MEMWBrd & IFIDrs2 != 5'h0 & _bypassAFromWB_T_5; // @[cpu.scala 328:50]
  wire  _bypassAFromMEM_T_2 = IFIDrs1 == EXMEMrd & _bypassAFromWB_T_1; // @[cpu.scala 330:29]
  wire [6:0] EXMEMop = io_rvfi_rst ? EXMEMIR[6:0] : EXMEMIR[6:0]; // @[cpu.scala 299:21 305:13 317:13]
  wire  _bypassAFromMEM_T_3 = EXMEMop == 7'h33; // @[cpu.scala 330:62]
  wire  bypassAFromMEM = IFIDrs1 == EXMEMrd & _bypassAFromWB_T_1 & EXMEMop == 7'h33; // @[cpu.scala 330:50]
  wire  _bypassBFromMEM_T_2 = IFIDrs2 == EXMEMrd & _bypassBFromWB_T_1; // @[cpu.scala 332:29]
  wire  bypassBFromMEM = IFIDrs2 == EXMEMrd & _bypassBFromWB_T_1 & _bypassAFromMEM_T_3; // @[cpu.scala 332:50]
  wire  _bypassAFromEX_T_2 = IFIDrs1 == IDEXrd & _bypassAFromWB_T_1; // @[cpu.scala 334:28]
  wire [6:0] IDEXop = io_rvfi_rst ? IDEXIR[6:0] : IDEXIR[6:0]; // @[cpu.scala 299:21 303:12 315:12]
  wire  _bypassAFromEX_T_3 = IDEXop == 7'h33; // @[cpu.scala 334:60]
  wire  bypassAFromEX = IFIDrs1 == IDEXrd & _bypassAFromWB_T_1 & IDEXop == 7'h33; // @[cpu.scala 334:49]
  wire  _bypassBFromEX_T_2 = IFIDrs2 == IDEXrd & _bypassBFromWB_T_1; // @[cpu.scala 336:28]
  wire  bypassBFromEX = IFIDrs2 == IDEXrd & _bypassBFromWB_T_1 & _bypassAFromEX_T_3; // @[cpu.scala 336:49]
  wire  _stall_T = EXMEMop == 7'h3; // @[cpu.scala 339:16]
  wire  _stall_T_8 = EXMEMop == 7'h3 & (_bypassAFromMEM_T_2 | _bypassBFromMEM_T_2); // @[cpu.scala 339:24]
  wire  _stall_T_9 = IDEXop == 7'h3; // @[cpu.scala 341:15]
  wire  _stall_T_17 = IDEXop == 7'h3 & (_bypassAFromEX_T_2 | _bypassBFromEX_T_2); // @[cpu.scala 341:23]
  wire  stall = _stall_T_8 | _stall_T_17; // @[cpu.scala 340:7]
  wire [6:0] IFIDop = io_rvfi_rst ? IFIDIR[6:0] : IFIDIR[6:0]; // @[cpu.scala 299:21 304:12 316:12]
  wire [63:0] _A_T_1 = IDEXA + IDEXB; // @[cpu.scala 382:20]
  wire [63:0] _GEN_5 = 5'h1 == IFIDrs1 ? Regs_1 : Regs_0; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_6 = 5'h2 == IFIDrs1 ? Regs_2 : _GEN_5; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_7 = 5'h3 == IFIDrs1 ? Regs_3 : _GEN_6; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_8 = 5'h4 == IFIDrs1 ? Regs_4 : _GEN_7; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_9 = 5'h5 == IFIDrs1 ? Regs_5 : _GEN_8; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_10 = 5'h6 == IFIDrs1 ? Regs_6 : _GEN_9; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_11 = 5'h7 == IFIDrs1 ? Regs_7 : _GEN_10; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_12 = 5'h8 == IFIDrs1 ? Regs_8 : _GEN_11; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_13 = 5'h9 == IFIDrs1 ? Regs_9 : _GEN_12; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_14 = 5'ha == IFIDrs1 ? Regs_10 : _GEN_13; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_15 = 5'hb == IFIDrs1 ? Regs_11 : _GEN_14; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_16 = 5'hc == IFIDrs1 ? Regs_12 : _GEN_15; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_17 = 5'hd == IFIDrs1 ? Regs_13 : _GEN_16; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_18 = 5'he == IFIDrs1 ? Regs_14 : _GEN_17; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_19 = 5'hf == IFIDrs1 ? Regs_15 : _GEN_18; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_20 = 5'h10 == IFIDrs1 ? Regs_16 : _GEN_19; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_21 = 5'h11 == IFIDrs1 ? Regs_17 : _GEN_20; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_22 = 5'h12 == IFIDrs1 ? Regs_18 : _GEN_21; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_23 = 5'h13 == IFIDrs1 ? Regs_19 : _GEN_22; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_24 = 5'h14 == IFIDrs1 ? Regs_20 : _GEN_23; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_25 = 5'h15 == IFIDrs1 ? Regs_21 : _GEN_24; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_26 = 5'h16 == IFIDrs1 ? Regs_22 : _GEN_25; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_27 = 5'h17 == IFIDrs1 ? Regs_23 : _GEN_26; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_28 = 5'h18 == IFIDrs1 ? Regs_24 : _GEN_27; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_29 = 5'h19 == IFIDrs1 ? Regs_25 : _GEN_28; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_30 = 5'h1a == IFIDrs1 ? Regs_26 : _GEN_29; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_31 = 5'h1b == IFIDrs1 ? Regs_27 : _GEN_30; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_32 = 5'h1c == IFIDrs1 ? Regs_28 : _GEN_31; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_33 = 5'h1d == IFIDrs1 ? Regs_29 : _GEN_32; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_34 = 5'h1e == IFIDrs1 ? Regs_30 : _GEN_33; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_35 = 5'h1f == IFIDrs1 ? Regs_31 : _GEN_34; // @[cpu.scala 390:{15,15}]
  wire [63:0] _GEN_37 = bypassAFromWB ? MEMWBValue : _GEN_35; // @[cpu.scala 386:33 388:11 391:11]
  wire [63:0] _GEN_39 = bypassAFromMEM ? EXMEMALUOut : _GEN_37; // @[cpu.scala 383:34 385:11]
  wire [63:0] _GEN_41 = bypassAFromEX ? _A_T_1 : _GEN_39; // @[cpu.scala 380:27 382:11]
  wire [63:0] A = ~stall ? _GEN_41 : 64'h0; // @[cpu.scala 353:27]
  wire [63:0] _B_T_1 = IDEXB + IDEXA; // @[cpu.scala 395:20]
  wire [63:0] _GEN_43 = 5'h1 == IFIDrs2 ? Regs_1 : Regs_0; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_44 = 5'h2 == IFIDrs2 ? Regs_2 : _GEN_43; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_45 = 5'h3 == IFIDrs2 ? Regs_3 : _GEN_44; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_46 = 5'h4 == IFIDrs2 ? Regs_4 : _GEN_45; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_47 = 5'h5 == IFIDrs2 ? Regs_5 : _GEN_46; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_48 = 5'h6 == IFIDrs2 ? Regs_6 : _GEN_47; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_49 = 5'h7 == IFIDrs2 ? Regs_7 : _GEN_48; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_50 = 5'h8 == IFIDrs2 ? Regs_8 : _GEN_49; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_51 = 5'h9 == IFIDrs2 ? Regs_9 : _GEN_50; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_52 = 5'ha == IFIDrs2 ? Regs_10 : _GEN_51; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_53 = 5'hb == IFIDrs2 ? Regs_11 : _GEN_52; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_54 = 5'hc == IFIDrs2 ? Regs_12 : _GEN_53; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_55 = 5'hd == IFIDrs2 ? Regs_13 : _GEN_54; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_56 = 5'he == IFIDrs2 ? Regs_14 : _GEN_55; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_57 = 5'hf == IFIDrs2 ? Regs_15 : _GEN_56; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_58 = 5'h10 == IFIDrs2 ? Regs_16 : _GEN_57; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_59 = 5'h11 == IFIDrs2 ? Regs_17 : _GEN_58; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_60 = 5'h12 == IFIDrs2 ? Regs_18 : _GEN_59; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_61 = 5'h13 == IFIDrs2 ? Regs_19 : _GEN_60; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_62 = 5'h14 == IFIDrs2 ? Regs_20 : _GEN_61; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_63 = 5'h15 == IFIDrs2 ? Regs_21 : _GEN_62; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_64 = 5'h16 == IFIDrs2 ? Regs_22 : _GEN_63; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_65 = 5'h17 == IFIDrs2 ? Regs_23 : _GEN_64; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_66 = 5'h18 == IFIDrs2 ? Regs_24 : _GEN_65; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_67 = 5'h19 == IFIDrs2 ? Regs_25 : _GEN_66; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_68 = 5'h1a == IFIDrs2 ? Regs_26 : _GEN_67; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_69 = 5'h1b == IFIDrs2 ? Regs_27 : _GEN_68; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_70 = 5'h1c == IFIDrs2 ? Regs_28 : _GEN_69; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_71 = 5'h1d == IFIDrs2 ? Regs_29 : _GEN_70; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_72 = 5'h1e == IFIDrs2 ? Regs_30 : _GEN_71; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_73 = 5'h1f == IFIDrs2 ? Regs_31 : _GEN_72; // @[cpu.scala 403:{15,15}]
  wire [63:0] _GEN_75 = bypassBFromWB ? MEMWBValue : _GEN_73; // @[cpu.scala 399:33 401:11 404:11]
  wire [63:0] _GEN_77 = bypassBFromMEM ? EXMEMALUOut : _GEN_75; // @[cpu.scala 396:34 398:11]
  wire [63:0] _GEN_79 = bypassBFromEX ? _B_T_1 : _GEN_77; // @[cpu.scala 393:27 395:11]
  wire [63:0] B = ~stall ? _GEN_79 : 64'h0; // @[cpu.scala 353:27]
  wire  takeBranch = IFIDop == 7'h63 & IFID_funct3 == 3'h0 & A == B; // @[cpu.scala 345:64]
  wire [12:0] _branchTarget_T_5 = {IFIDIR[31],1'h0,IFIDIR[30:25],IFIDIR[11:7]}; // @[cpu.scala 367:11]
  wire [63:0] _GEN_6363 = {{51{_branchTarget_T_5[12]}},_branchTarget_T_5}; // @[cpu.scala 362:42]
  wire [63:0] branchTarget = $signed(CurPC) + $signed(_GEN_6363); // @[cpu.scala 367:19]
  wire [11:0] _EXMEMALUOut_T_2 = IDEXIR[31:20]; // @[cpu.scala 415:53]
  wire [63:0] _GEN_6364 = {{52{_EXMEMALUOut_T_2[11]}},_EXMEMALUOut_T_2}; // @[cpu.scala 415:36]
  wire [63:0] _EXMEMALUOut_T_6 = $signed(IDEXA) + $signed(_GEN_6364); // @[cpu.scala 415:61]
  wire [11:0] _EXMEMALUOut_T_11 = {IDEXIR[31:25],IDEXrd}; // @[cpu.scala 420:9]
  wire [63:0] _GEN_6365 = {{52{_EXMEMALUOut_T_11[11]}},_EXMEMALUOut_T_11}; // @[cpu.scala 417:36]
  wire [63:0] _EXMEMALUOut_T_15 = $signed(IDEXA) + $signed(_GEN_6365); // @[cpu.scala 420:17]
  wire [31:0] _GEN_94 = 10'h1 == EXMEMALUOut[9:0] ? DMemory_1 : DMemory_0; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_95 = 10'h2 == EXMEMALUOut[9:0] ? DMemory_2 : _GEN_94; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_96 = 10'h3 == EXMEMALUOut[9:0] ? DMemory_3 : _GEN_95; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_97 = 10'h4 == EXMEMALUOut[9:0] ? DMemory_4 : _GEN_96; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_98 = 10'h5 == EXMEMALUOut[9:0] ? DMemory_5 : _GEN_97; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_99 = 10'h6 == EXMEMALUOut[9:0] ? DMemory_6 : _GEN_98; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_100 = 10'h7 == EXMEMALUOut[9:0] ? DMemory_7 : _GEN_99; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_101 = 10'h8 == EXMEMALUOut[9:0] ? DMemory_8 : _GEN_100; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_102 = 10'h9 == EXMEMALUOut[9:0] ? DMemory_9 : _GEN_101; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_103 = 10'ha == EXMEMALUOut[9:0] ? DMemory_10 : _GEN_102; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_104 = 10'hb == EXMEMALUOut[9:0] ? DMemory_11 : _GEN_103; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_105 = 10'hc == EXMEMALUOut[9:0] ? DMemory_12 : _GEN_104; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_106 = 10'hd == EXMEMALUOut[9:0] ? DMemory_13 : _GEN_105; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_107 = 10'he == EXMEMALUOut[9:0] ? DMemory_14 : _GEN_106; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_108 = 10'hf == EXMEMALUOut[9:0] ? DMemory_15 : _GEN_107; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_109 = 10'h10 == EXMEMALUOut[9:0] ? DMemory_16 : _GEN_108; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_110 = 10'h11 == EXMEMALUOut[9:0] ? DMemory_17 : _GEN_109; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_111 = 10'h12 == EXMEMALUOut[9:0] ? DMemory_18 : _GEN_110; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_112 = 10'h13 == EXMEMALUOut[9:0] ? DMemory_19 : _GEN_111; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_113 = 10'h14 == EXMEMALUOut[9:0] ? DMemory_20 : _GEN_112; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_114 = 10'h15 == EXMEMALUOut[9:0] ? DMemory_21 : _GEN_113; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_115 = 10'h16 == EXMEMALUOut[9:0] ? DMemory_22 : _GEN_114; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_116 = 10'h17 == EXMEMALUOut[9:0] ? DMemory_23 : _GEN_115; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_117 = 10'h18 == EXMEMALUOut[9:0] ? DMemory_24 : _GEN_116; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_118 = 10'h19 == EXMEMALUOut[9:0] ? DMemory_25 : _GEN_117; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_119 = 10'h1a == EXMEMALUOut[9:0] ? DMemory_26 : _GEN_118; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_120 = 10'h1b == EXMEMALUOut[9:0] ? DMemory_27 : _GEN_119; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_121 = 10'h1c == EXMEMALUOut[9:0] ? DMemory_28 : _GEN_120; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_122 = 10'h1d == EXMEMALUOut[9:0] ? DMemory_29 : _GEN_121; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_123 = 10'h1e == EXMEMALUOut[9:0] ? DMemory_30 : _GEN_122; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_124 = 10'h1f == EXMEMALUOut[9:0] ? DMemory_31 : _GEN_123; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_125 = 10'h20 == EXMEMALUOut[9:0] ? DMemory_32 : _GEN_124; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_126 = 10'h21 == EXMEMALUOut[9:0] ? DMemory_33 : _GEN_125; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_127 = 10'h22 == EXMEMALUOut[9:0] ? DMemory_34 : _GEN_126; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_128 = 10'h23 == EXMEMALUOut[9:0] ? DMemory_35 : _GEN_127; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_129 = 10'h24 == EXMEMALUOut[9:0] ? DMemory_36 : _GEN_128; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_130 = 10'h25 == EXMEMALUOut[9:0] ? DMemory_37 : _GEN_129; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_131 = 10'h26 == EXMEMALUOut[9:0] ? DMemory_38 : _GEN_130; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_132 = 10'h27 == EXMEMALUOut[9:0] ? DMemory_39 : _GEN_131; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_133 = 10'h28 == EXMEMALUOut[9:0] ? DMemory_40 : _GEN_132; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_134 = 10'h29 == EXMEMALUOut[9:0] ? DMemory_41 : _GEN_133; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_135 = 10'h2a == EXMEMALUOut[9:0] ? DMemory_42 : _GEN_134; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_136 = 10'h2b == EXMEMALUOut[9:0] ? DMemory_43 : _GEN_135; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_137 = 10'h2c == EXMEMALUOut[9:0] ? DMemory_44 : _GEN_136; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_138 = 10'h2d == EXMEMALUOut[9:0] ? DMemory_45 : _GEN_137; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_139 = 10'h2e == EXMEMALUOut[9:0] ? DMemory_46 : _GEN_138; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_140 = 10'h2f == EXMEMALUOut[9:0] ? DMemory_47 : _GEN_139; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_141 = 10'h30 == EXMEMALUOut[9:0] ? DMemory_48 : _GEN_140; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_142 = 10'h31 == EXMEMALUOut[9:0] ? DMemory_49 : _GEN_141; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_143 = 10'h32 == EXMEMALUOut[9:0] ? DMemory_50 : _GEN_142; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_144 = 10'h33 == EXMEMALUOut[9:0] ? DMemory_51 : _GEN_143; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_145 = 10'h34 == EXMEMALUOut[9:0] ? DMemory_52 : _GEN_144; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_146 = 10'h35 == EXMEMALUOut[9:0] ? DMemory_53 : _GEN_145; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_147 = 10'h36 == EXMEMALUOut[9:0] ? DMemory_54 : _GEN_146; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_148 = 10'h37 == EXMEMALUOut[9:0] ? DMemory_55 : _GEN_147; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_149 = 10'h38 == EXMEMALUOut[9:0] ? DMemory_56 : _GEN_148; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_150 = 10'h39 == EXMEMALUOut[9:0] ? DMemory_57 : _GEN_149; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_151 = 10'h3a == EXMEMALUOut[9:0] ? DMemory_58 : _GEN_150; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_152 = 10'h3b == EXMEMALUOut[9:0] ? DMemory_59 : _GEN_151; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_153 = 10'h3c == EXMEMALUOut[9:0] ? DMemory_60 : _GEN_152; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_154 = 10'h3d == EXMEMALUOut[9:0] ? DMemory_61 : _GEN_153; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_155 = 10'h3e == EXMEMALUOut[9:0] ? DMemory_62 : _GEN_154; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_156 = 10'h3f == EXMEMALUOut[9:0] ? DMemory_63 : _GEN_155; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_157 = 10'h40 == EXMEMALUOut[9:0] ? DMemory_64 : _GEN_156; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_158 = 10'h41 == EXMEMALUOut[9:0] ? DMemory_65 : _GEN_157; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_159 = 10'h42 == EXMEMALUOut[9:0] ? DMemory_66 : _GEN_158; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_160 = 10'h43 == EXMEMALUOut[9:0] ? DMemory_67 : _GEN_159; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_161 = 10'h44 == EXMEMALUOut[9:0] ? DMemory_68 : _GEN_160; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_162 = 10'h45 == EXMEMALUOut[9:0] ? DMemory_69 : _GEN_161; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_163 = 10'h46 == EXMEMALUOut[9:0] ? DMemory_70 : _GEN_162; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_164 = 10'h47 == EXMEMALUOut[9:0] ? DMemory_71 : _GEN_163; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_165 = 10'h48 == EXMEMALUOut[9:0] ? DMemory_72 : _GEN_164; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_166 = 10'h49 == EXMEMALUOut[9:0] ? DMemory_73 : _GEN_165; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_167 = 10'h4a == EXMEMALUOut[9:0] ? DMemory_74 : _GEN_166; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_168 = 10'h4b == EXMEMALUOut[9:0] ? DMemory_75 : _GEN_167; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_169 = 10'h4c == EXMEMALUOut[9:0] ? DMemory_76 : _GEN_168; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_170 = 10'h4d == EXMEMALUOut[9:0] ? DMemory_77 : _GEN_169; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_171 = 10'h4e == EXMEMALUOut[9:0] ? DMemory_78 : _GEN_170; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_172 = 10'h4f == EXMEMALUOut[9:0] ? DMemory_79 : _GEN_171; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_173 = 10'h50 == EXMEMALUOut[9:0] ? DMemory_80 : _GEN_172; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_174 = 10'h51 == EXMEMALUOut[9:0] ? DMemory_81 : _GEN_173; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_175 = 10'h52 == EXMEMALUOut[9:0] ? DMemory_82 : _GEN_174; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_176 = 10'h53 == EXMEMALUOut[9:0] ? DMemory_83 : _GEN_175; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_177 = 10'h54 == EXMEMALUOut[9:0] ? DMemory_84 : _GEN_176; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_178 = 10'h55 == EXMEMALUOut[9:0] ? DMemory_85 : _GEN_177; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_179 = 10'h56 == EXMEMALUOut[9:0] ? DMemory_86 : _GEN_178; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_180 = 10'h57 == EXMEMALUOut[9:0] ? DMemory_87 : _GEN_179; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_181 = 10'h58 == EXMEMALUOut[9:0] ? DMemory_88 : _GEN_180; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_182 = 10'h59 == EXMEMALUOut[9:0] ? DMemory_89 : _GEN_181; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_183 = 10'h5a == EXMEMALUOut[9:0] ? DMemory_90 : _GEN_182; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_184 = 10'h5b == EXMEMALUOut[9:0] ? DMemory_91 : _GEN_183; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_185 = 10'h5c == EXMEMALUOut[9:0] ? DMemory_92 : _GEN_184; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_186 = 10'h5d == EXMEMALUOut[9:0] ? DMemory_93 : _GEN_185; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_187 = 10'h5e == EXMEMALUOut[9:0] ? DMemory_94 : _GEN_186; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_188 = 10'h5f == EXMEMALUOut[9:0] ? DMemory_95 : _GEN_187; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_189 = 10'h60 == EXMEMALUOut[9:0] ? DMemory_96 : _GEN_188; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_190 = 10'h61 == EXMEMALUOut[9:0] ? DMemory_97 : _GEN_189; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_191 = 10'h62 == EXMEMALUOut[9:0] ? DMemory_98 : _GEN_190; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_192 = 10'h63 == EXMEMALUOut[9:0] ? DMemory_99 : _GEN_191; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_193 = 10'h64 == EXMEMALUOut[9:0] ? DMemory_100 : _GEN_192; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_194 = 10'h65 == EXMEMALUOut[9:0] ? DMemory_101 : _GEN_193; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_195 = 10'h66 == EXMEMALUOut[9:0] ? DMemory_102 : _GEN_194; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_196 = 10'h67 == EXMEMALUOut[9:0] ? DMemory_103 : _GEN_195; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_197 = 10'h68 == EXMEMALUOut[9:0] ? DMemory_104 : _GEN_196; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_198 = 10'h69 == EXMEMALUOut[9:0] ? DMemory_105 : _GEN_197; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_199 = 10'h6a == EXMEMALUOut[9:0] ? DMemory_106 : _GEN_198; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_200 = 10'h6b == EXMEMALUOut[9:0] ? DMemory_107 : _GEN_199; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_201 = 10'h6c == EXMEMALUOut[9:0] ? DMemory_108 : _GEN_200; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_202 = 10'h6d == EXMEMALUOut[9:0] ? DMemory_109 : _GEN_201; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_203 = 10'h6e == EXMEMALUOut[9:0] ? DMemory_110 : _GEN_202; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_204 = 10'h6f == EXMEMALUOut[9:0] ? DMemory_111 : _GEN_203; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_205 = 10'h70 == EXMEMALUOut[9:0] ? DMemory_112 : _GEN_204; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_206 = 10'h71 == EXMEMALUOut[9:0] ? DMemory_113 : _GEN_205; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_207 = 10'h72 == EXMEMALUOut[9:0] ? DMemory_114 : _GEN_206; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_208 = 10'h73 == EXMEMALUOut[9:0] ? DMemory_115 : _GEN_207; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_209 = 10'h74 == EXMEMALUOut[9:0] ? DMemory_116 : _GEN_208; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_210 = 10'h75 == EXMEMALUOut[9:0] ? DMemory_117 : _GEN_209; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_211 = 10'h76 == EXMEMALUOut[9:0] ? DMemory_118 : _GEN_210; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_212 = 10'h77 == EXMEMALUOut[9:0] ? DMemory_119 : _GEN_211; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_213 = 10'h78 == EXMEMALUOut[9:0] ? DMemory_120 : _GEN_212; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_214 = 10'h79 == EXMEMALUOut[9:0] ? DMemory_121 : _GEN_213; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_215 = 10'h7a == EXMEMALUOut[9:0] ? DMemory_122 : _GEN_214; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_216 = 10'h7b == EXMEMALUOut[9:0] ? DMemory_123 : _GEN_215; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_217 = 10'h7c == EXMEMALUOut[9:0] ? DMemory_124 : _GEN_216; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_218 = 10'h7d == EXMEMALUOut[9:0] ? DMemory_125 : _GEN_217; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_219 = 10'h7e == EXMEMALUOut[9:0] ? DMemory_126 : _GEN_218; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_220 = 10'h7f == EXMEMALUOut[9:0] ? DMemory_127 : _GEN_219; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_221 = 10'h80 == EXMEMALUOut[9:0] ? DMemory_128 : _GEN_220; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_222 = 10'h81 == EXMEMALUOut[9:0] ? DMemory_129 : _GEN_221; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_223 = 10'h82 == EXMEMALUOut[9:0] ? DMemory_130 : _GEN_222; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_224 = 10'h83 == EXMEMALUOut[9:0] ? DMemory_131 : _GEN_223; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_225 = 10'h84 == EXMEMALUOut[9:0] ? DMemory_132 : _GEN_224; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_226 = 10'h85 == EXMEMALUOut[9:0] ? DMemory_133 : _GEN_225; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_227 = 10'h86 == EXMEMALUOut[9:0] ? DMemory_134 : _GEN_226; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_228 = 10'h87 == EXMEMALUOut[9:0] ? DMemory_135 : _GEN_227; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_229 = 10'h88 == EXMEMALUOut[9:0] ? DMemory_136 : _GEN_228; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_230 = 10'h89 == EXMEMALUOut[9:0] ? DMemory_137 : _GEN_229; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_231 = 10'h8a == EXMEMALUOut[9:0] ? DMemory_138 : _GEN_230; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_232 = 10'h8b == EXMEMALUOut[9:0] ? DMemory_139 : _GEN_231; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_233 = 10'h8c == EXMEMALUOut[9:0] ? DMemory_140 : _GEN_232; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_234 = 10'h8d == EXMEMALUOut[9:0] ? DMemory_141 : _GEN_233; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_235 = 10'h8e == EXMEMALUOut[9:0] ? DMemory_142 : _GEN_234; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_236 = 10'h8f == EXMEMALUOut[9:0] ? DMemory_143 : _GEN_235; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_237 = 10'h90 == EXMEMALUOut[9:0] ? DMemory_144 : _GEN_236; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_238 = 10'h91 == EXMEMALUOut[9:0] ? DMemory_145 : _GEN_237; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_239 = 10'h92 == EXMEMALUOut[9:0] ? DMemory_146 : _GEN_238; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_240 = 10'h93 == EXMEMALUOut[9:0] ? DMemory_147 : _GEN_239; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_241 = 10'h94 == EXMEMALUOut[9:0] ? DMemory_148 : _GEN_240; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_242 = 10'h95 == EXMEMALUOut[9:0] ? DMemory_149 : _GEN_241; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_243 = 10'h96 == EXMEMALUOut[9:0] ? DMemory_150 : _GEN_242; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_244 = 10'h97 == EXMEMALUOut[9:0] ? DMemory_151 : _GEN_243; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_245 = 10'h98 == EXMEMALUOut[9:0] ? DMemory_152 : _GEN_244; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_246 = 10'h99 == EXMEMALUOut[9:0] ? DMemory_153 : _GEN_245; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_247 = 10'h9a == EXMEMALUOut[9:0] ? DMemory_154 : _GEN_246; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_248 = 10'h9b == EXMEMALUOut[9:0] ? DMemory_155 : _GEN_247; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_249 = 10'h9c == EXMEMALUOut[9:0] ? DMemory_156 : _GEN_248; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_250 = 10'h9d == EXMEMALUOut[9:0] ? DMemory_157 : _GEN_249; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_251 = 10'h9e == EXMEMALUOut[9:0] ? DMemory_158 : _GEN_250; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_252 = 10'h9f == EXMEMALUOut[9:0] ? DMemory_159 : _GEN_251; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_253 = 10'ha0 == EXMEMALUOut[9:0] ? DMemory_160 : _GEN_252; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_254 = 10'ha1 == EXMEMALUOut[9:0] ? DMemory_161 : _GEN_253; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_255 = 10'ha2 == EXMEMALUOut[9:0] ? DMemory_162 : _GEN_254; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_256 = 10'ha3 == EXMEMALUOut[9:0] ? DMemory_163 : _GEN_255; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_257 = 10'ha4 == EXMEMALUOut[9:0] ? DMemory_164 : _GEN_256; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_258 = 10'ha5 == EXMEMALUOut[9:0] ? DMemory_165 : _GEN_257; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_259 = 10'ha6 == EXMEMALUOut[9:0] ? DMemory_166 : _GEN_258; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_260 = 10'ha7 == EXMEMALUOut[9:0] ? DMemory_167 : _GEN_259; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_261 = 10'ha8 == EXMEMALUOut[9:0] ? DMemory_168 : _GEN_260; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_262 = 10'ha9 == EXMEMALUOut[9:0] ? DMemory_169 : _GEN_261; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_263 = 10'haa == EXMEMALUOut[9:0] ? DMemory_170 : _GEN_262; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_264 = 10'hab == EXMEMALUOut[9:0] ? DMemory_171 : _GEN_263; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_265 = 10'hac == EXMEMALUOut[9:0] ? DMemory_172 : _GEN_264; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_266 = 10'had == EXMEMALUOut[9:0] ? DMemory_173 : _GEN_265; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_267 = 10'hae == EXMEMALUOut[9:0] ? DMemory_174 : _GEN_266; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_268 = 10'haf == EXMEMALUOut[9:0] ? DMemory_175 : _GEN_267; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_269 = 10'hb0 == EXMEMALUOut[9:0] ? DMemory_176 : _GEN_268; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_270 = 10'hb1 == EXMEMALUOut[9:0] ? DMemory_177 : _GEN_269; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_271 = 10'hb2 == EXMEMALUOut[9:0] ? DMemory_178 : _GEN_270; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_272 = 10'hb3 == EXMEMALUOut[9:0] ? DMemory_179 : _GEN_271; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_273 = 10'hb4 == EXMEMALUOut[9:0] ? DMemory_180 : _GEN_272; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_274 = 10'hb5 == EXMEMALUOut[9:0] ? DMemory_181 : _GEN_273; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_275 = 10'hb6 == EXMEMALUOut[9:0] ? DMemory_182 : _GEN_274; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_276 = 10'hb7 == EXMEMALUOut[9:0] ? DMemory_183 : _GEN_275; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_277 = 10'hb8 == EXMEMALUOut[9:0] ? DMemory_184 : _GEN_276; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_278 = 10'hb9 == EXMEMALUOut[9:0] ? DMemory_185 : _GEN_277; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_279 = 10'hba == EXMEMALUOut[9:0] ? DMemory_186 : _GEN_278; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_280 = 10'hbb == EXMEMALUOut[9:0] ? DMemory_187 : _GEN_279; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_281 = 10'hbc == EXMEMALUOut[9:0] ? DMemory_188 : _GEN_280; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_282 = 10'hbd == EXMEMALUOut[9:0] ? DMemory_189 : _GEN_281; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_283 = 10'hbe == EXMEMALUOut[9:0] ? DMemory_190 : _GEN_282; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_284 = 10'hbf == EXMEMALUOut[9:0] ? DMemory_191 : _GEN_283; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_285 = 10'hc0 == EXMEMALUOut[9:0] ? DMemory_192 : _GEN_284; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_286 = 10'hc1 == EXMEMALUOut[9:0] ? DMemory_193 : _GEN_285; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_287 = 10'hc2 == EXMEMALUOut[9:0] ? DMemory_194 : _GEN_286; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_288 = 10'hc3 == EXMEMALUOut[9:0] ? DMemory_195 : _GEN_287; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_289 = 10'hc4 == EXMEMALUOut[9:0] ? DMemory_196 : _GEN_288; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_290 = 10'hc5 == EXMEMALUOut[9:0] ? DMemory_197 : _GEN_289; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_291 = 10'hc6 == EXMEMALUOut[9:0] ? DMemory_198 : _GEN_290; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_292 = 10'hc7 == EXMEMALUOut[9:0] ? DMemory_199 : _GEN_291; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_293 = 10'hc8 == EXMEMALUOut[9:0] ? DMemory_200 : _GEN_292; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_294 = 10'hc9 == EXMEMALUOut[9:0] ? DMemory_201 : _GEN_293; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_295 = 10'hca == EXMEMALUOut[9:0] ? DMemory_202 : _GEN_294; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_296 = 10'hcb == EXMEMALUOut[9:0] ? DMemory_203 : _GEN_295; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_297 = 10'hcc == EXMEMALUOut[9:0] ? DMemory_204 : _GEN_296; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_298 = 10'hcd == EXMEMALUOut[9:0] ? DMemory_205 : _GEN_297; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_299 = 10'hce == EXMEMALUOut[9:0] ? DMemory_206 : _GEN_298; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_300 = 10'hcf == EXMEMALUOut[9:0] ? DMemory_207 : _GEN_299; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_301 = 10'hd0 == EXMEMALUOut[9:0] ? DMemory_208 : _GEN_300; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_302 = 10'hd1 == EXMEMALUOut[9:0] ? DMemory_209 : _GEN_301; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_303 = 10'hd2 == EXMEMALUOut[9:0] ? DMemory_210 : _GEN_302; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_304 = 10'hd3 == EXMEMALUOut[9:0] ? DMemory_211 : _GEN_303; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_305 = 10'hd4 == EXMEMALUOut[9:0] ? DMemory_212 : _GEN_304; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_306 = 10'hd5 == EXMEMALUOut[9:0] ? DMemory_213 : _GEN_305; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_307 = 10'hd6 == EXMEMALUOut[9:0] ? DMemory_214 : _GEN_306; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_308 = 10'hd7 == EXMEMALUOut[9:0] ? DMemory_215 : _GEN_307; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_309 = 10'hd8 == EXMEMALUOut[9:0] ? DMemory_216 : _GEN_308; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_310 = 10'hd9 == EXMEMALUOut[9:0] ? DMemory_217 : _GEN_309; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_311 = 10'hda == EXMEMALUOut[9:0] ? DMemory_218 : _GEN_310; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_312 = 10'hdb == EXMEMALUOut[9:0] ? DMemory_219 : _GEN_311; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_313 = 10'hdc == EXMEMALUOut[9:0] ? DMemory_220 : _GEN_312; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_314 = 10'hdd == EXMEMALUOut[9:0] ? DMemory_221 : _GEN_313; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_315 = 10'hde == EXMEMALUOut[9:0] ? DMemory_222 : _GEN_314; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_316 = 10'hdf == EXMEMALUOut[9:0] ? DMemory_223 : _GEN_315; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_317 = 10'he0 == EXMEMALUOut[9:0] ? DMemory_224 : _GEN_316; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_318 = 10'he1 == EXMEMALUOut[9:0] ? DMemory_225 : _GEN_317; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_319 = 10'he2 == EXMEMALUOut[9:0] ? DMemory_226 : _GEN_318; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_320 = 10'he3 == EXMEMALUOut[9:0] ? DMemory_227 : _GEN_319; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_321 = 10'he4 == EXMEMALUOut[9:0] ? DMemory_228 : _GEN_320; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_322 = 10'he5 == EXMEMALUOut[9:0] ? DMemory_229 : _GEN_321; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_323 = 10'he6 == EXMEMALUOut[9:0] ? DMemory_230 : _GEN_322; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_324 = 10'he7 == EXMEMALUOut[9:0] ? DMemory_231 : _GEN_323; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_325 = 10'he8 == EXMEMALUOut[9:0] ? DMemory_232 : _GEN_324; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_326 = 10'he9 == EXMEMALUOut[9:0] ? DMemory_233 : _GEN_325; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_327 = 10'hea == EXMEMALUOut[9:0] ? DMemory_234 : _GEN_326; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_328 = 10'heb == EXMEMALUOut[9:0] ? DMemory_235 : _GEN_327; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_329 = 10'hec == EXMEMALUOut[9:0] ? DMemory_236 : _GEN_328; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_330 = 10'hed == EXMEMALUOut[9:0] ? DMemory_237 : _GEN_329; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_331 = 10'hee == EXMEMALUOut[9:0] ? DMemory_238 : _GEN_330; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_332 = 10'hef == EXMEMALUOut[9:0] ? DMemory_239 : _GEN_331; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_333 = 10'hf0 == EXMEMALUOut[9:0] ? DMemory_240 : _GEN_332; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_334 = 10'hf1 == EXMEMALUOut[9:0] ? DMemory_241 : _GEN_333; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_335 = 10'hf2 == EXMEMALUOut[9:0] ? DMemory_242 : _GEN_334; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_336 = 10'hf3 == EXMEMALUOut[9:0] ? DMemory_243 : _GEN_335; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_337 = 10'hf4 == EXMEMALUOut[9:0] ? DMemory_244 : _GEN_336; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_338 = 10'hf5 == EXMEMALUOut[9:0] ? DMemory_245 : _GEN_337; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_339 = 10'hf6 == EXMEMALUOut[9:0] ? DMemory_246 : _GEN_338; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_340 = 10'hf7 == EXMEMALUOut[9:0] ? DMemory_247 : _GEN_339; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_341 = 10'hf8 == EXMEMALUOut[9:0] ? DMemory_248 : _GEN_340; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_342 = 10'hf9 == EXMEMALUOut[9:0] ? DMemory_249 : _GEN_341; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_343 = 10'hfa == EXMEMALUOut[9:0] ? DMemory_250 : _GEN_342; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_344 = 10'hfb == EXMEMALUOut[9:0] ? DMemory_251 : _GEN_343; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_345 = 10'hfc == EXMEMALUOut[9:0] ? DMemory_252 : _GEN_344; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_346 = 10'hfd == EXMEMALUOut[9:0] ? DMemory_253 : _GEN_345; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_347 = 10'hfe == EXMEMALUOut[9:0] ? DMemory_254 : _GEN_346; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_348 = 10'hff == EXMEMALUOut[9:0] ? DMemory_255 : _GEN_347; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_349 = 10'h100 == EXMEMALUOut[9:0] ? DMemory_256 : _GEN_348; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_350 = 10'h101 == EXMEMALUOut[9:0] ? DMemory_257 : _GEN_349; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_351 = 10'h102 == EXMEMALUOut[9:0] ? DMemory_258 : _GEN_350; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_352 = 10'h103 == EXMEMALUOut[9:0] ? DMemory_259 : _GEN_351; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_353 = 10'h104 == EXMEMALUOut[9:0] ? DMemory_260 : _GEN_352; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_354 = 10'h105 == EXMEMALUOut[9:0] ? DMemory_261 : _GEN_353; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_355 = 10'h106 == EXMEMALUOut[9:0] ? DMemory_262 : _GEN_354; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_356 = 10'h107 == EXMEMALUOut[9:0] ? DMemory_263 : _GEN_355; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_357 = 10'h108 == EXMEMALUOut[9:0] ? DMemory_264 : _GEN_356; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_358 = 10'h109 == EXMEMALUOut[9:0] ? DMemory_265 : _GEN_357; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_359 = 10'h10a == EXMEMALUOut[9:0] ? DMemory_266 : _GEN_358; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_360 = 10'h10b == EXMEMALUOut[9:0] ? DMemory_267 : _GEN_359; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_361 = 10'h10c == EXMEMALUOut[9:0] ? DMemory_268 : _GEN_360; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_362 = 10'h10d == EXMEMALUOut[9:0] ? DMemory_269 : _GEN_361; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_363 = 10'h10e == EXMEMALUOut[9:0] ? DMemory_270 : _GEN_362; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_364 = 10'h10f == EXMEMALUOut[9:0] ? DMemory_271 : _GEN_363; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_365 = 10'h110 == EXMEMALUOut[9:0] ? DMemory_272 : _GEN_364; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_366 = 10'h111 == EXMEMALUOut[9:0] ? DMemory_273 : _GEN_365; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_367 = 10'h112 == EXMEMALUOut[9:0] ? DMemory_274 : _GEN_366; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_368 = 10'h113 == EXMEMALUOut[9:0] ? DMemory_275 : _GEN_367; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_369 = 10'h114 == EXMEMALUOut[9:0] ? DMemory_276 : _GEN_368; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_370 = 10'h115 == EXMEMALUOut[9:0] ? DMemory_277 : _GEN_369; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_371 = 10'h116 == EXMEMALUOut[9:0] ? DMemory_278 : _GEN_370; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_372 = 10'h117 == EXMEMALUOut[9:0] ? DMemory_279 : _GEN_371; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_373 = 10'h118 == EXMEMALUOut[9:0] ? DMemory_280 : _GEN_372; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_374 = 10'h119 == EXMEMALUOut[9:0] ? DMemory_281 : _GEN_373; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_375 = 10'h11a == EXMEMALUOut[9:0] ? DMemory_282 : _GEN_374; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_376 = 10'h11b == EXMEMALUOut[9:0] ? DMemory_283 : _GEN_375; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_377 = 10'h11c == EXMEMALUOut[9:0] ? DMemory_284 : _GEN_376; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_378 = 10'h11d == EXMEMALUOut[9:0] ? DMemory_285 : _GEN_377; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_379 = 10'h11e == EXMEMALUOut[9:0] ? DMemory_286 : _GEN_378; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_380 = 10'h11f == EXMEMALUOut[9:0] ? DMemory_287 : _GEN_379; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_381 = 10'h120 == EXMEMALUOut[9:0] ? DMemory_288 : _GEN_380; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_382 = 10'h121 == EXMEMALUOut[9:0] ? DMemory_289 : _GEN_381; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_383 = 10'h122 == EXMEMALUOut[9:0] ? DMemory_290 : _GEN_382; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_384 = 10'h123 == EXMEMALUOut[9:0] ? DMemory_291 : _GEN_383; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_385 = 10'h124 == EXMEMALUOut[9:0] ? DMemory_292 : _GEN_384; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_386 = 10'h125 == EXMEMALUOut[9:0] ? DMemory_293 : _GEN_385; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_387 = 10'h126 == EXMEMALUOut[9:0] ? DMemory_294 : _GEN_386; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_388 = 10'h127 == EXMEMALUOut[9:0] ? DMemory_295 : _GEN_387; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_389 = 10'h128 == EXMEMALUOut[9:0] ? DMemory_296 : _GEN_388; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_390 = 10'h129 == EXMEMALUOut[9:0] ? DMemory_297 : _GEN_389; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_391 = 10'h12a == EXMEMALUOut[9:0] ? DMemory_298 : _GEN_390; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_392 = 10'h12b == EXMEMALUOut[9:0] ? DMemory_299 : _GEN_391; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_393 = 10'h12c == EXMEMALUOut[9:0] ? DMemory_300 : _GEN_392; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_394 = 10'h12d == EXMEMALUOut[9:0] ? DMemory_301 : _GEN_393; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_395 = 10'h12e == EXMEMALUOut[9:0] ? DMemory_302 : _GEN_394; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_396 = 10'h12f == EXMEMALUOut[9:0] ? DMemory_303 : _GEN_395; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_397 = 10'h130 == EXMEMALUOut[9:0] ? DMemory_304 : _GEN_396; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_398 = 10'h131 == EXMEMALUOut[9:0] ? DMemory_305 : _GEN_397; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_399 = 10'h132 == EXMEMALUOut[9:0] ? DMemory_306 : _GEN_398; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_400 = 10'h133 == EXMEMALUOut[9:0] ? DMemory_307 : _GEN_399; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_401 = 10'h134 == EXMEMALUOut[9:0] ? DMemory_308 : _GEN_400; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_402 = 10'h135 == EXMEMALUOut[9:0] ? DMemory_309 : _GEN_401; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_403 = 10'h136 == EXMEMALUOut[9:0] ? DMemory_310 : _GEN_402; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_404 = 10'h137 == EXMEMALUOut[9:0] ? DMemory_311 : _GEN_403; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_405 = 10'h138 == EXMEMALUOut[9:0] ? DMemory_312 : _GEN_404; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_406 = 10'h139 == EXMEMALUOut[9:0] ? DMemory_313 : _GEN_405; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_407 = 10'h13a == EXMEMALUOut[9:0] ? DMemory_314 : _GEN_406; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_408 = 10'h13b == EXMEMALUOut[9:0] ? DMemory_315 : _GEN_407; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_409 = 10'h13c == EXMEMALUOut[9:0] ? DMemory_316 : _GEN_408; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_410 = 10'h13d == EXMEMALUOut[9:0] ? DMemory_317 : _GEN_409; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_411 = 10'h13e == EXMEMALUOut[9:0] ? DMemory_318 : _GEN_410; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_412 = 10'h13f == EXMEMALUOut[9:0] ? DMemory_319 : _GEN_411; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_413 = 10'h140 == EXMEMALUOut[9:0] ? DMemory_320 : _GEN_412; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_414 = 10'h141 == EXMEMALUOut[9:0] ? DMemory_321 : _GEN_413; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_415 = 10'h142 == EXMEMALUOut[9:0] ? DMemory_322 : _GEN_414; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_416 = 10'h143 == EXMEMALUOut[9:0] ? DMemory_323 : _GEN_415; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_417 = 10'h144 == EXMEMALUOut[9:0] ? DMemory_324 : _GEN_416; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_418 = 10'h145 == EXMEMALUOut[9:0] ? DMemory_325 : _GEN_417; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_419 = 10'h146 == EXMEMALUOut[9:0] ? DMemory_326 : _GEN_418; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_420 = 10'h147 == EXMEMALUOut[9:0] ? DMemory_327 : _GEN_419; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_421 = 10'h148 == EXMEMALUOut[9:0] ? DMemory_328 : _GEN_420; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_422 = 10'h149 == EXMEMALUOut[9:0] ? DMemory_329 : _GEN_421; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_423 = 10'h14a == EXMEMALUOut[9:0] ? DMemory_330 : _GEN_422; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_424 = 10'h14b == EXMEMALUOut[9:0] ? DMemory_331 : _GEN_423; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_425 = 10'h14c == EXMEMALUOut[9:0] ? DMemory_332 : _GEN_424; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_426 = 10'h14d == EXMEMALUOut[9:0] ? DMemory_333 : _GEN_425; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_427 = 10'h14e == EXMEMALUOut[9:0] ? DMemory_334 : _GEN_426; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_428 = 10'h14f == EXMEMALUOut[9:0] ? DMemory_335 : _GEN_427; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_429 = 10'h150 == EXMEMALUOut[9:0] ? DMemory_336 : _GEN_428; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_430 = 10'h151 == EXMEMALUOut[9:0] ? DMemory_337 : _GEN_429; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_431 = 10'h152 == EXMEMALUOut[9:0] ? DMemory_338 : _GEN_430; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_432 = 10'h153 == EXMEMALUOut[9:0] ? DMemory_339 : _GEN_431; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_433 = 10'h154 == EXMEMALUOut[9:0] ? DMemory_340 : _GEN_432; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_434 = 10'h155 == EXMEMALUOut[9:0] ? DMemory_341 : _GEN_433; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_435 = 10'h156 == EXMEMALUOut[9:0] ? DMemory_342 : _GEN_434; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_436 = 10'h157 == EXMEMALUOut[9:0] ? DMemory_343 : _GEN_435; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_437 = 10'h158 == EXMEMALUOut[9:0] ? DMemory_344 : _GEN_436; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_438 = 10'h159 == EXMEMALUOut[9:0] ? DMemory_345 : _GEN_437; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_439 = 10'h15a == EXMEMALUOut[9:0] ? DMemory_346 : _GEN_438; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_440 = 10'h15b == EXMEMALUOut[9:0] ? DMemory_347 : _GEN_439; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_441 = 10'h15c == EXMEMALUOut[9:0] ? DMemory_348 : _GEN_440; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_442 = 10'h15d == EXMEMALUOut[9:0] ? DMemory_349 : _GEN_441; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_443 = 10'h15e == EXMEMALUOut[9:0] ? DMemory_350 : _GEN_442; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_444 = 10'h15f == EXMEMALUOut[9:0] ? DMemory_351 : _GEN_443; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_445 = 10'h160 == EXMEMALUOut[9:0] ? DMemory_352 : _GEN_444; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_446 = 10'h161 == EXMEMALUOut[9:0] ? DMemory_353 : _GEN_445; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_447 = 10'h162 == EXMEMALUOut[9:0] ? DMemory_354 : _GEN_446; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_448 = 10'h163 == EXMEMALUOut[9:0] ? DMemory_355 : _GEN_447; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_449 = 10'h164 == EXMEMALUOut[9:0] ? DMemory_356 : _GEN_448; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_450 = 10'h165 == EXMEMALUOut[9:0] ? DMemory_357 : _GEN_449; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_451 = 10'h166 == EXMEMALUOut[9:0] ? DMemory_358 : _GEN_450; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_452 = 10'h167 == EXMEMALUOut[9:0] ? DMemory_359 : _GEN_451; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_453 = 10'h168 == EXMEMALUOut[9:0] ? DMemory_360 : _GEN_452; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_454 = 10'h169 == EXMEMALUOut[9:0] ? DMemory_361 : _GEN_453; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_455 = 10'h16a == EXMEMALUOut[9:0] ? DMemory_362 : _GEN_454; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_456 = 10'h16b == EXMEMALUOut[9:0] ? DMemory_363 : _GEN_455; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_457 = 10'h16c == EXMEMALUOut[9:0] ? DMemory_364 : _GEN_456; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_458 = 10'h16d == EXMEMALUOut[9:0] ? DMemory_365 : _GEN_457; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_459 = 10'h16e == EXMEMALUOut[9:0] ? DMemory_366 : _GEN_458; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_460 = 10'h16f == EXMEMALUOut[9:0] ? DMemory_367 : _GEN_459; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_461 = 10'h170 == EXMEMALUOut[9:0] ? DMemory_368 : _GEN_460; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_462 = 10'h171 == EXMEMALUOut[9:0] ? DMemory_369 : _GEN_461; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_463 = 10'h172 == EXMEMALUOut[9:0] ? DMemory_370 : _GEN_462; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_464 = 10'h173 == EXMEMALUOut[9:0] ? DMemory_371 : _GEN_463; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_465 = 10'h174 == EXMEMALUOut[9:0] ? DMemory_372 : _GEN_464; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_466 = 10'h175 == EXMEMALUOut[9:0] ? DMemory_373 : _GEN_465; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_467 = 10'h176 == EXMEMALUOut[9:0] ? DMemory_374 : _GEN_466; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_468 = 10'h177 == EXMEMALUOut[9:0] ? DMemory_375 : _GEN_467; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_469 = 10'h178 == EXMEMALUOut[9:0] ? DMemory_376 : _GEN_468; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_470 = 10'h179 == EXMEMALUOut[9:0] ? DMemory_377 : _GEN_469; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_471 = 10'h17a == EXMEMALUOut[9:0] ? DMemory_378 : _GEN_470; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_472 = 10'h17b == EXMEMALUOut[9:0] ? DMemory_379 : _GEN_471; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_473 = 10'h17c == EXMEMALUOut[9:0] ? DMemory_380 : _GEN_472; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_474 = 10'h17d == EXMEMALUOut[9:0] ? DMemory_381 : _GEN_473; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_475 = 10'h17e == EXMEMALUOut[9:0] ? DMemory_382 : _GEN_474; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_476 = 10'h17f == EXMEMALUOut[9:0] ? DMemory_383 : _GEN_475; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_477 = 10'h180 == EXMEMALUOut[9:0] ? DMemory_384 : _GEN_476; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_478 = 10'h181 == EXMEMALUOut[9:0] ? DMemory_385 : _GEN_477; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_479 = 10'h182 == EXMEMALUOut[9:0] ? DMemory_386 : _GEN_478; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_480 = 10'h183 == EXMEMALUOut[9:0] ? DMemory_387 : _GEN_479; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_481 = 10'h184 == EXMEMALUOut[9:0] ? DMemory_388 : _GEN_480; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_482 = 10'h185 == EXMEMALUOut[9:0] ? DMemory_389 : _GEN_481; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_483 = 10'h186 == EXMEMALUOut[9:0] ? DMemory_390 : _GEN_482; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_484 = 10'h187 == EXMEMALUOut[9:0] ? DMemory_391 : _GEN_483; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_485 = 10'h188 == EXMEMALUOut[9:0] ? DMemory_392 : _GEN_484; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_486 = 10'h189 == EXMEMALUOut[9:0] ? DMemory_393 : _GEN_485; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_487 = 10'h18a == EXMEMALUOut[9:0] ? DMemory_394 : _GEN_486; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_488 = 10'h18b == EXMEMALUOut[9:0] ? DMemory_395 : _GEN_487; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_489 = 10'h18c == EXMEMALUOut[9:0] ? DMemory_396 : _GEN_488; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_490 = 10'h18d == EXMEMALUOut[9:0] ? DMemory_397 : _GEN_489; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_491 = 10'h18e == EXMEMALUOut[9:0] ? DMemory_398 : _GEN_490; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_492 = 10'h18f == EXMEMALUOut[9:0] ? DMemory_399 : _GEN_491; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_493 = 10'h190 == EXMEMALUOut[9:0] ? DMemory_400 : _GEN_492; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_494 = 10'h191 == EXMEMALUOut[9:0] ? DMemory_401 : _GEN_493; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_495 = 10'h192 == EXMEMALUOut[9:0] ? DMemory_402 : _GEN_494; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_496 = 10'h193 == EXMEMALUOut[9:0] ? DMemory_403 : _GEN_495; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_497 = 10'h194 == EXMEMALUOut[9:0] ? DMemory_404 : _GEN_496; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_498 = 10'h195 == EXMEMALUOut[9:0] ? DMemory_405 : _GEN_497; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_499 = 10'h196 == EXMEMALUOut[9:0] ? DMemory_406 : _GEN_498; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_500 = 10'h197 == EXMEMALUOut[9:0] ? DMemory_407 : _GEN_499; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_501 = 10'h198 == EXMEMALUOut[9:0] ? DMemory_408 : _GEN_500; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_502 = 10'h199 == EXMEMALUOut[9:0] ? DMemory_409 : _GEN_501; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_503 = 10'h19a == EXMEMALUOut[9:0] ? DMemory_410 : _GEN_502; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_504 = 10'h19b == EXMEMALUOut[9:0] ? DMemory_411 : _GEN_503; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_505 = 10'h19c == EXMEMALUOut[9:0] ? DMemory_412 : _GEN_504; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_506 = 10'h19d == EXMEMALUOut[9:0] ? DMemory_413 : _GEN_505; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_507 = 10'h19e == EXMEMALUOut[9:0] ? DMemory_414 : _GEN_506; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_508 = 10'h19f == EXMEMALUOut[9:0] ? DMemory_415 : _GEN_507; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_509 = 10'h1a0 == EXMEMALUOut[9:0] ? DMemory_416 : _GEN_508; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_510 = 10'h1a1 == EXMEMALUOut[9:0] ? DMemory_417 : _GEN_509; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_511 = 10'h1a2 == EXMEMALUOut[9:0] ? DMemory_418 : _GEN_510; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_512 = 10'h1a3 == EXMEMALUOut[9:0] ? DMemory_419 : _GEN_511; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_513 = 10'h1a4 == EXMEMALUOut[9:0] ? DMemory_420 : _GEN_512; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_514 = 10'h1a5 == EXMEMALUOut[9:0] ? DMemory_421 : _GEN_513; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_515 = 10'h1a6 == EXMEMALUOut[9:0] ? DMemory_422 : _GEN_514; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_516 = 10'h1a7 == EXMEMALUOut[9:0] ? DMemory_423 : _GEN_515; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_517 = 10'h1a8 == EXMEMALUOut[9:0] ? DMemory_424 : _GEN_516; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_518 = 10'h1a9 == EXMEMALUOut[9:0] ? DMemory_425 : _GEN_517; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_519 = 10'h1aa == EXMEMALUOut[9:0] ? DMemory_426 : _GEN_518; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_520 = 10'h1ab == EXMEMALUOut[9:0] ? DMemory_427 : _GEN_519; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_521 = 10'h1ac == EXMEMALUOut[9:0] ? DMemory_428 : _GEN_520; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_522 = 10'h1ad == EXMEMALUOut[9:0] ? DMemory_429 : _GEN_521; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_523 = 10'h1ae == EXMEMALUOut[9:0] ? DMemory_430 : _GEN_522; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_524 = 10'h1af == EXMEMALUOut[9:0] ? DMemory_431 : _GEN_523; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_525 = 10'h1b0 == EXMEMALUOut[9:0] ? DMemory_432 : _GEN_524; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_526 = 10'h1b1 == EXMEMALUOut[9:0] ? DMemory_433 : _GEN_525; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_527 = 10'h1b2 == EXMEMALUOut[9:0] ? DMemory_434 : _GEN_526; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_528 = 10'h1b3 == EXMEMALUOut[9:0] ? DMemory_435 : _GEN_527; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_529 = 10'h1b4 == EXMEMALUOut[9:0] ? DMemory_436 : _GEN_528; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_530 = 10'h1b5 == EXMEMALUOut[9:0] ? DMemory_437 : _GEN_529; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_531 = 10'h1b6 == EXMEMALUOut[9:0] ? DMemory_438 : _GEN_530; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_532 = 10'h1b7 == EXMEMALUOut[9:0] ? DMemory_439 : _GEN_531; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_533 = 10'h1b8 == EXMEMALUOut[9:0] ? DMemory_440 : _GEN_532; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_534 = 10'h1b9 == EXMEMALUOut[9:0] ? DMemory_441 : _GEN_533; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_535 = 10'h1ba == EXMEMALUOut[9:0] ? DMemory_442 : _GEN_534; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_536 = 10'h1bb == EXMEMALUOut[9:0] ? DMemory_443 : _GEN_535; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_537 = 10'h1bc == EXMEMALUOut[9:0] ? DMemory_444 : _GEN_536; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_538 = 10'h1bd == EXMEMALUOut[9:0] ? DMemory_445 : _GEN_537; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_539 = 10'h1be == EXMEMALUOut[9:0] ? DMemory_446 : _GEN_538; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_540 = 10'h1bf == EXMEMALUOut[9:0] ? DMemory_447 : _GEN_539; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_541 = 10'h1c0 == EXMEMALUOut[9:0] ? DMemory_448 : _GEN_540; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_542 = 10'h1c1 == EXMEMALUOut[9:0] ? DMemory_449 : _GEN_541; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_543 = 10'h1c2 == EXMEMALUOut[9:0] ? DMemory_450 : _GEN_542; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_544 = 10'h1c3 == EXMEMALUOut[9:0] ? DMemory_451 : _GEN_543; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_545 = 10'h1c4 == EXMEMALUOut[9:0] ? DMemory_452 : _GEN_544; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_546 = 10'h1c5 == EXMEMALUOut[9:0] ? DMemory_453 : _GEN_545; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_547 = 10'h1c6 == EXMEMALUOut[9:0] ? DMemory_454 : _GEN_546; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_548 = 10'h1c7 == EXMEMALUOut[9:0] ? DMemory_455 : _GEN_547; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_549 = 10'h1c8 == EXMEMALUOut[9:0] ? DMemory_456 : _GEN_548; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_550 = 10'h1c9 == EXMEMALUOut[9:0] ? DMemory_457 : _GEN_549; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_551 = 10'h1ca == EXMEMALUOut[9:0] ? DMemory_458 : _GEN_550; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_552 = 10'h1cb == EXMEMALUOut[9:0] ? DMemory_459 : _GEN_551; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_553 = 10'h1cc == EXMEMALUOut[9:0] ? DMemory_460 : _GEN_552; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_554 = 10'h1cd == EXMEMALUOut[9:0] ? DMemory_461 : _GEN_553; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_555 = 10'h1ce == EXMEMALUOut[9:0] ? DMemory_462 : _GEN_554; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_556 = 10'h1cf == EXMEMALUOut[9:0] ? DMemory_463 : _GEN_555; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_557 = 10'h1d0 == EXMEMALUOut[9:0] ? DMemory_464 : _GEN_556; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_558 = 10'h1d1 == EXMEMALUOut[9:0] ? DMemory_465 : _GEN_557; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_559 = 10'h1d2 == EXMEMALUOut[9:0] ? DMemory_466 : _GEN_558; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_560 = 10'h1d3 == EXMEMALUOut[9:0] ? DMemory_467 : _GEN_559; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_561 = 10'h1d4 == EXMEMALUOut[9:0] ? DMemory_468 : _GEN_560; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_562 = 10'h1d5 == EXMEMALUOut[9:0] ? DMemory_469 : _GEN_561; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_563 = 10'h1d6 == EXMEMALUOut[9:0] ? DMemory_470 : _GEN_562; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_564 = 10'h1d7 == EXMEMALUOut[9:0] ? DMemory_471 : _GEN_563; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_565 = 10'h1d8 == EXMEMALUOut[9:0] ? DMemory_472 : _GEN_564; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_566 = 10'h1d9 == EXMEMALUOut[9:0] ? DMemory_473 : _GEN_565; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_567 = 10'h1da == EXMEMALUOut[9:0] ? DMemory_474 : _GEN_566; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_568 = 10'h1db == EXMEMALUOut[9:0] ? DMemory_475 : _GEN_567; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_569 = 10'h1dc == EXMEMALUOut[9:0] ? DMemory_476 : _GEN_568; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_570 = 10'h1dd == EXMEMALUOut[9:0] ? DMemory_477 : _GEN_569; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_571 = 10'h1de == EXMEMALUOut[9:0] ? DMemory_478 : _GEN_570; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_572 = 10'h1df == EXMEMALUOut[9:0] ? DMemory_479 : _GEN_571; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_573 = 10'h1e0 == EXMEMALUOut[9:0] ? DMemory_480 : _GEN_572; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_574 = 10'h1e1 == EXMEMALUOut[9:0] ? DMemory_481 : _GEN_573; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_575 = 10'h1e2 == EXMEMALUOut[9:0] ? DMemory_482 : _GEN_574; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_576 = 10'h1e3 == EXMEMALUOut[9:0] ? DMemory_483 : _GEN_575; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_577 = 10'h1e4 == EXMEMALUOut[9:0] ? DMemory_484 : _GEN_576; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_578 = 10'h1e5 == EXMEMALUOut[9:0] ? DMemory_485 : _GEN_577; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_579 = 10'h1e6 == EXMEMALUOut[9:0] ? DMemory_486 : _GEN_578; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_580 = 10'h1e7 == EXMEMALUOut[9:0] ? DMemory_487 : _GEN_579; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_581 = 10'h1e8 == EXMEMALUOut[9:0] ? DMemory_488 : _GEN_580; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_582 = 10'h1e9 == EXMEMALUOut[9:0] ? DMemory_489 : _GEN_581; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_583 = 10'h1ea == EXMEMALUOut[9:0] ? DMemory_490 : _GEN_582; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_584 = 10'h1eb == EXMEMALUOut[9:0] ? DMemory_491 : _GEN_583; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_585 = 10'h1ec == EXMEMALUOut[9:0] ? DMemory_492 : _GEN_584; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_586 = 10'h1ed == EXMEMALUOut[9:0] ? DMemory_493 : _GEN_585; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_587 = 10'h1ee == EXMEMALUOut[9:0] ? DMemory_494 : _GEN_586; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_588 = 10'h1ef == EXMEMALUOut[9:0] ? DMemory_495 : _GEN_587; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_589 = 10'h1f0 == EXMEMALUOut[9:0] ? DMemory_496 : _GEN_588; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_590 = 10'h1f1 == EXMEMALUOut[9:0] ? DMemory_497 : _GEN_589; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_591 = 10'h1f2 == EXMEMALUOut[9:0] ? DMemory_498 : _GEN_590; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_592 = 10'h1f3 == EXMEMALUOut[9:0] ? DMemory_499 : _GEN_591; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_593 = 10'h1f4 == EXMEMALUOut[9:0] ? DMemory_500 : _GEN_592; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_594 = 10'h1f5 == EXMEMALUOut[9:0] ? DMemory_501 : _GEN_593; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_595 = 10'h1f6 == EXMEMALUOut[9:0] ? DMemory_502 : _GEN_594; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_596 = 10'h1f7 == EXMEMALUOut[9:0] ? DMemory_503 : _GEN_595; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_597 = 10'h1f8 == EXMEMALUOut[9:0] ? DMemory_504 : _GEN_596; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_598 = 10'h1f9 == EXMEMALUOut[9:0] ? DMemory_505 : _GEN_597; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_599 = 10'h1fa == EXMEMALUOut[9:0] ? DMemory_506 : _GEN_598; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_600 = 10'h1fb == EXMEMALUOut[9:0] ? DMemory_507 : _GEN_599; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_601 = 10'h1fc == EXMEMALUOut[9:0] ? DMemory_508 : _GEN_600; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_602 = 10'h1fd == EXMEMALUOut[9:0] ? DMemory_509 : _GEN_601; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_603 = 10'h1fe == EXMEMALUOut[9:0] ? DMemory_510 : _GEN_602; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_604 = 10'h1ff == EXMEMALUOut[9:0] ? DMemory_511 : _GEN_603; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_605 = 10'h200 == EXMEMALUOut[9:0] ? DMemory_512 : _GEN_604; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_606 = 10'h201 == EXMEMALUOut[9:0] ? DMemory_513 : _GEN_605; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_607 = 10'h202 == EXMEMALUOut[9:0] ? DMemory_514 : _GEN_606; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_608 = 10'h203 == EXMEMALUOut[9:0] ? DMemory_515 : _GEN_607; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_609 = 10'h204 == EXMEMALUOut[9:0] ? DMemory_516 : _GEN_608; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_610 = 10'h205 == EXMEMALUOut[9:0] ? DMemory_517 : _GEN_609; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_611 = 10'h206 == EXMEMALUOut[9:0] ? DMemory_518 : _GEN_610; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_612 = 10'h207 == EXMEMALUOut[9:0] ? DMemory_519 : _GEN_611; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_613 = 10'h208 == EXMEMALUOut[9:0] ? DMemory_520 : _GEN_612; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_614 = 10'h209 == EXMEMALUOut[9:0] ? DMemory_521 : _GEN_613; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_615 = 10'h20a == EXMEMALUOut[9:0] ? DMemory_522 : _GEN_614; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_616 = 10'h20b == EXMEMALUOut[9:0] ? DMemory_523 : _GEN_615; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_617 = 10'h20c == EXMEMALUOut[9:0] ? DMemory_524 : _GEN_616; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_618 = 10'h20d == EXMEMALUOut[9:0] ? DMemory_525 : _GEN_617; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_619 = 10'h20e == EXMEMALUOut[9:0] ? DMemory_526 : _GEN_618; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_620 = 10'h20f == EXMEMALUOut[9:0] ? DMemory_527 : _GEN_619; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_621 = 10'h210 == EXMEMALUOut[9:0] ? DMemory_528 : _GEN_620; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_622 = 10'h211 == EXMEMALUOut[9:0] ? DMemory_529 : _GEN_621; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_623 = 10'h212 == EXMEMALUOut[9:0] ? DMemory_530 : _GEN_622; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_624 = 10'h213 == EXMEMALUOut[9:0] ? DMemory_531 : _GEN_623; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_625 = 10'h214 == EXMEMALUOut[9:0] ? DMemory_532 : _GEN_624; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_626 = 10'h215 == EXMEMALUOut[9:0] ? DMemory_533 : _GEN_625; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_627 = 10'h216 == EXMEMALUOut[9:0] ? DMemory_534 : _GEN_626; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_628 = 10'h217 == EXMEMALUOut[9:0] ? DMemory_535 : _GEN_627; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_629 = 10'h218 == EXMEMALUOut[9:0] ? DMemory_536 : _GEN_628; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_630 = 10'h219 == EXMEMALUOut[9:0] ? DMemory_537 : _GEN_629; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_631 = 10'h21a == EXMEMALUOut[9:0] ? DMemory_538 : _GEN_630; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_632 = 10'h21b == EXMEMALUOut[9:0] ? DMemory_539 : _GEN_631; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_633 = 10'h21c == EXMEMALUOut[9:0] ? DMemory_540 : _GEN_632; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_634 = 10'h21d == EXMEMALUOut[9:0] ? DMemory_541 : _GEN_633; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_635 = 10'h21e == EXMEMALUOut[9:0] ? DMemory_542 : _GEN_634; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_636 = 10'h21f == EXMEMALUOut[9:0] ? DMemory_543 : _GEN_635; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_637 = 10'h220 == EXMEMALUOut[9:0] ? DMemory_544 : _GEN_636; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_638 = 10'h221 == EXMEMALUOut[9:0] ? DMemory_545 : _GEN_637; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_639 = 10'h222 == EXMEMALUOut[9:0] ? DMemory_546 : _GEN_638; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_640 = 10'h223 == EXMEMALUOut[9:0] ? DMemory_547 : _GEN_639; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_641 = 10'h224 == EXMEMALUOut[9:0] ? DMemory_548 : _GEN_640; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_642 = 10'h225 == EXMEMALUOut[9:0] ? DMemory_549 : _GEN_641; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_643 = 10'h226 == EXMEMALUOut[9:0] ? DMemory_550 : _GEN_642; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_644 = 10'h227 == EXMEMALUOut[9:0] ? DMemory_551 : _GEN_643; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_645 = 10'h228 == EXMEMALUOut[9:0] ? DMemory_552 : _GEN_644; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_646 = 10'h229 == EXMEMALUOut[9:0] ? DMemory_553 : _GEN_645; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_647 = 10'h22a == EXMEMALUOut[9:0] ? DMemory_554 : _GEN_646; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_648 = 10'h22b == EXMEMALUOut[9:0] ? DMemory_555 : _GEN_647; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_649 = 10'h22c == EXMEMALUOut[9:0] ? DMemory_556 : _GEN_648; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_650 = 10'h22d == EXMEMALUOut[9:0] ? DMemory_557 : _GEN_649; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_651 = 10'h22e == EXMEMALUOut[9:0] ? DMemory_558 : _GEN_650; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_652 = 10'h22f == EXMEMALUOut[9:0] ? DMemory_559 : _GEN_651; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_653 = 10'h230 == EXMEMALUOut[9:0] ? DMemory_560 : _GEN_652; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_654 = 10'h231 == EXMEMALUOut[9:0] ? DMemory_561 : _GEN_653; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_655 = 10'h232 == EXMEMALUOut[9:0] ? DMemory_562 : _GEN_654; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_656 = 10'h233 == EXMEMALUOut[9:0] ? DMemory_563 : _GEN_655; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_657 = 10'h234 == EXMEMALUOut[9:0] ? DMemory_564 : _GEN_656; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_658 = 10'h235 == EXMEMALUOut[9:0] ? DMemory_565 : _GEN_657; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_659 = 10'h236 == EXMEMALUOut[9:0] ? DMemory_566 : _GEN_658; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_660 = 10'h237 == EXMEMALUOut[9:0] ? DMemory_567 : _GEN_659; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_661 = 10'h238 == EXMEMALUOut[9:0] ? DMemory_568 : _GEN_660; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_662 = 10'h239 == EXMEMALUOut[9:0] ? DMemory_569 : _GEN_661; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_663 = 10'h23a == EXMEMALUOut[9:0] ? DMemory_570 : _GEN_662; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_664 = 10'h23b == EXMEMALUOut[9:0] ? DMemory_571 : _GEN_663; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_665 = 10'h23c == EXMEMALUOut[9:0] ? DMemory_572 : _GEN_664; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_666 = 10'h23d == EXMEMALUOut[9:0] ? DMemory_573 : _GEN_665; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_667 = 10'h23e == EXMEMALUOut[9:0] ? DMemory_574 : _GEN_666; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_668 = 10'h23f == EXMEMALUOut[9:0] ? DMemory_575 : _GEN_667; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_669 = 10'h240 == EXMEMALUOut[9:0] ? DMemory_576 : _GEN_668; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_670 = 10'h241 == EXMEMALUOut[9:0] ? DMemory_577 : _GEN_669; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_671 = 10'h242 == EXMEMALUOut[9:0] ? DMemory_578 : _GEN_670; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_672 = 10'h243 == EXMEMALUOut[9:0] ? DMemory_579 : _GEN_671; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_673 = 10'h244 == EXMEMALUOut[9:0] ? DMemory_580 : _GEN_672; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_674 = 10'h245 == EXMEMALUOut[9:0] ? DMemory_581 : _GEN_673; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_675 = 10'h246 == EXMEMALUOut[9:0] ? DMemory_582 : _GEN_674; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_676 = 10'h247 == EXMEMALUOut[9:0] ? DMemory_583 : _GEN_675; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_677 = 10'h248 == EXMEMALUOut[9:0] ? DMemory_584 : _GEN_676; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_678 = 10'h249 == EXMEMALUOut[9:0] ? DMemory_585 : _GEN_677; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_679 = 10'h24a == EXMEMALUOut[9:0] ? DMemory_586 : _GEN_678; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_680 = 10'h24b == EXMEMALUOut[9:0] ? DMemory_587 : _GEN_679; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_681 = 10'h24c == EXMEMALUOut[9:0] ? DMemory_588 : _GEN_680; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_682 = 10'h24d == EXMEMALUOut[9:0] ? DMemory_589 : _GEN_681; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_683 = 10'h24e == EXMEMALUOut[9:0] ? DMemory_590 : _GEN_682; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_684 = 10'h24f == EXMEMALUOut[9:0] ? DMemory_591 : _GEN_683; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_685 = 10'h250 == EXMEMALUOut[9:0] ? DMemory_592 : _GEN_684; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_686 = 10'h251 == EXMEMALUOut[9:0] ? DMemory_593 : _GEN_685; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_687 = 10'h252 == EXMEMALUOut[9:0] ? DMemory_594 : _GEN_686; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_688 = 10'h253 == EXMEMALUOut[9:0] ? DMemory_595 : _GEN_687; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_689 = 10'h254 == EXMEMALUOut[9:0] ? DMemory_596 : _GEN_688; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_690 = 10'h255 == EXMEMALUOut[9:0] ? DMemory_597 : _GEN_689; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_691 = 10'h256 == EXMEMALUOut[9:0] ? DMemory_598 : _GEN_690; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_692 = 10'h257 == EXMEMALUOut[9:0] ? DMemory_599 : _GEN_691; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_693 = 10'h258 == EXMEMALUOut[9:0] ? DMemory_600 : _GEN_692; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_694 = 10'h259 == EXMEMALUOut[9:0] ? DMemory_601 : _GEN_693; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_695 = 10'h25a == EXMEMALUOut[9:0] ? DMemory_602 : _GEN_694; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_696 = 10'h25b == EXMEMALUOut[9:0] ? DMemory_603 : _GEN_695; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_697 = 10'h25c == EXMEMALUOut[9:0] ? DMemory_604 : _GEN_696; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_698 = 10'h25d == EXMEMALUOut[9:0] ? DMemory_605 : _GEN_697; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_699 = 10'h25e == EXMEMALUOut[9:0] ? DMemory_606 : _GEN_698; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_700 = 10'h25f == EXMEMALUOut[9:0] ? DMemory_607 : _GEN_699; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_701 = 10'h260 == EXMEMALUOut[9:0] ? DMemory_608 : _GEN_700; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_702 = 10'h261 == EXMEMALUOut[9:0] ? DMemory_609 : _GEN_701; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_703 = 10'h262 == EXMEMALUOut[9:0] ? DMemory_610 : _GEN_702; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_704 = 10'h263 == EXMEMALUOut[9:0] ? DMemory_611 : _GEN_703; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_705 = 10'h264 == EXMEMALUOut[9:0] ? DMemory_612 : _GEN_704; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_706 = 10'h265 == EXMEMALUOut[9:0] ? DMemory_613 : _GEN_705; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_707 = 10'h266 == EXMEMALUOut[9:0] ? DMemory_614 : _GEN_706; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_708 = 10'h267 == EXMEMALUOut[9:0] ? DMemory_615 : _GEN_707; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_709 = 10'h268 == EXMEMALUOut[9:0] ? DMemory_616 : _GEN_708; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_710 = 10'h269 == EXMEMALUOut[9:0] ? DMemory_617 : _GEN_709; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_711 = 10'h26a == EXMEMALUOut[9:0] ? DMemory_618 : _GEN_710; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_712 = 10'h26b == EXMEMALUOut[9:0] ? DMemory_619 : _GEN_711; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_713 = 10'h26c == EXMEMALUOut[9:0] ? DMemory_620 : _GEN_712; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_714 = 10'h26d == EXMEMALUOut[9:0] ? DMemory_621 : _GEN_713; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_715 = 10'h26e == EXMEMALUOut[9:0] ? DMemory_622 : _GEN_714; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_716 = 10'h26f == EXMEMALUOut[9:0] ? DMemory_623 : _GEN_715; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_717 = 10'h270 == EXMEMALUOut[9:0] ? DMemory_624 : _GEN_716; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_718 = 10'h271 == EXMEMALUOut[9:0] ? DMemory_625 : _GEN_717; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_719 = 10'h272 == EXMEMALUOut[9:0] ? DMemory_626 : _GEN_718; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_720 = 10'h273 == EXMEMALUOut[9:0] ? DMemory_627 : _GEN_719; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_721 = 10'h274 == EXMEMALUOut[9:0] ? DMemory_628 : _GEN_720; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_722 = 10'h275 == EXMEMALUOut[9:0] ? DMemory_629 : _GEN_721; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_723 = 10'h276 == EXMEMALUOut[9:0] ? DMemory_630 : _GEN_722; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_724 = 10'h277 == EXMEMALUOut[9:0] ? DMemory_631 : _GEN_723; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_725 = 10'h278 == EXMEMALUOut[9:0] ? DMemory_632 : _GEN_724; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_726 = 10'h279 == EXMEMALUOut[9:0] ? DMemory_633 : _GEN_725; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_727 = 10'h27a == EXMEMALUOut[9:0] ? DMemory_634 : _GEN_726; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_728 = 10'h27b == EXMEMALUOut[9:0] ? DMemory_635 : _GEN_727; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_729 = 10'h27c == EXMEMALUOut[9:0] ? DMemory_636 : _GEN_728; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_730 = 10'h27d == EXMEMALUOut[9:0] ? DMemory_637 : _GEN_729; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_731 = 10'h27e == EXMEMALUOut[9:0] ? DMemory_638 : _GEN_730; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_732 = 10'h27f == EXMEMALUOut[9:0] ? DMemory_639 : _GEN_731; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_733 = 10'h280 == EXMEMALUOut[9:0] ? DMemory_640 : _GEN_732; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_734 = 10'h281 == EXMEMALUOut[9:0] ? DMemory_641 : _GEN_733; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_735 = 10'h282 == EXMEMALUOut[9:0] ? DMemory_642 : _GEN_734; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_736 = 10'h283 == EXMEMALUOut[9:0] ? DMemory_643 : _GEN_735; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_737 = 10'h284 == EXMEMALUOut[9:0] ? DMemory_644 : _GEN_736; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_738 = 10'h285 == EXMEMALUOut[9:0] ? DMemory_645 : _GEN_737; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_739 = 10'h286 == EXMEMALUOut[9:0] ? DMemory_646 : _GEN_738; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_740 = 10'h287 == EXMEMALUOut[9:0] ? DMemory_647 : _GEN_739; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_741 = 10'h288 == EXMEMALUOut[9:0] ? DMemory_648 : _GEN_740; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_742 = 10'h289 == EXMEMALUOut[9:0] ? DMemory_649 : _GEN_741; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_743 = 10'h28a == EXMEMALUOut[9:0] ? DMemory_650 : _GEN_742; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_744 = 10'h28b == EXMEMALUOut[9:0] ? DMemory_651 : _GEN_743; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_745 = 10'h28c == EXMEMALUOut[9:0] ? DMemory_652 : _GEN_744; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_746 = 10'h28d == EXMEMALUOut[9:0] ? DMemory_653 : _GEN_745; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_747 = 10'h28e == EXMEMALUOut[9:0] ? DMemory_654 : _GEN_746; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_748 = 10'h28f == EXMEMALUOut[9:0] ? DMemory_655 : _GEN_747; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_749 = 10'h290 == EXMEMALUOut[9:0] ? DMemory_656 : _GEN_748; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_750 = 10'h291 == EXMEMALUOut[9:0] ? DMemory_657 : _GEN_749; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_751 = 10'h292 == EXMEMALUOut[9:0] ? DMemory_658 : _GEN_750; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_752 = 10'h293 == EXMEMALUOut[9:0] ? DMemory_659 : _GEN_751; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_753 = 10'h294 == EXMEMALUOut[9:0] ? DMemory_660 : _GEN_752; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_754 = 10'h295 == EXMEMALUOut[9:0] ? DMemory_661 : _GEN_753; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_755 = 10'h296 == EXMEMALUOut[9:0] ? DMemory_662 : _GEN_754; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_756 = 10'h297 == EXMEMALUOut[9:0] ? DMemory_663 : _GEN_755; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_757 = 10'h298 == EXMEMALUOut[9:0] ? DMemory_664 : _GEN_756; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_758 = 10'h299 == EXMEMALUOut[9:0] ? DMemory_665 : _GEN_757; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_759 = 10'h29a == EXMEMALUOut[9:0] ? DMemory_666 : _GEN_758; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_760 = 10'h29b == EXMEMALUOut[9:0] ? DMemory_667 : _GEN_759; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_761 = 10'h29c == EXMEMALUOut[9:0] ? DMemory_668 : _GEN_760; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_762 = 10'h29d == EXMEMALUOut[9:0] ? DMemory_669 : _GEN_761; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_763 = 10'h29e == EXMEMALUOut[9:0] ? DMemory_670 : _GEN_762; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_764 = 10'h29f == EXMEMALUOut[9:0] ? DMemory_671 : _GEN_763; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_765 = 10'h2a0 == EXMEMALUOut[9:0] ? DMemory_672 : _GEN_764; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_766 = 10'h2a1 == EXMEMALUOut[9:0] ? DMemory_673 : _GEN_765; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_767 = 10'h2a2 == EXMEMALUOut[9:0] ? DMemory_674 : _GEN_766; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_768 = 10'h2a3 == EXMEMALUOut[9:0] ? DMemory_675 : _GEN_767; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_769 = 10'h2a4 == EXMEMALUOut[9:0] ? DMemory_676 : _GEN_768; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_770 = 10'h2a5 == EXMEMALUOut[9:0] ? DMemory_677 : _GEN_769; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_771 = 10'h2a6 == EXMEMALUOut[9:0] ? DMemory_678 : _GEN_770; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_772 = 10'h2a7 == EXMEMALUOut[9:0] ? DMemory_679 : _GEN_771; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_773 = 10'h2a8 == EXMEMALUOut[9:0] ? DMemory_680 : _GEN_772; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_774 = 10'h2a9 == EXMEMALUOut[9:0] ? DMemory_681 : _GEN_773; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_775 = 10'h2aa == EXMEMALUOut[9:0] ? DMemory_682 : _GEN_774; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_776 = 10'h2ab == EXMEMALUOut[9:0] ? DMemory_683 : _GEN_775; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_777 = 10'h2ac == EXMEMALUOut[9:0] ? DMemory_684 : _GEN_776; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_778 = 10'h2ad == EXMEMALUOut[9:0] ? DMemory_685 : _GEN_777; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_779 = 10'h2ae == EXMEMALUOut[9:0] ? DMemory_686 : _GEN_778; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_780 = 10'h2af == EXMEMALUOut[9:0] ? DMemory_687 : _GEN_779; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_781 = 10'h2b0 == EXMEMALUOut[9:0] ? DMemory_688 : _GEN_780; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_782 = 10'h2b1 == EXMEMALUOut[9:0] ? DMemory_689 : _GEN_781; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_783 = 10'h2b2 == EXMEMALUOut[9:0] ? DMemory_690 : _GEN_782; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_784 = 10'h2b3 == EXMEMALUOut[9:0] ? DMemory_691 : _GEN_783; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_785 = 10'h2b4 == EXMEMALUOut[9:0] ? DMemory_692 : _GEN_784; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_786 = 10'h2b5 == EXMEMALUOut[9:0] ? DMemory_693 : _GEN_785; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_787 = 10'h2b6 == EXMEMALUOut[9:0] ? DMemory_694 : _GEN_786; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_788 = 10'h2b7 == EXMEMALUOut[9:0] ? DMemory_695 : _GEN_787; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_789 = 10'h2b8 == EXMEMALUOut[9:0] ? DMemory_696 : _GEN_788; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_790 = 10'h2b9 == EXMEMALUOut[9:0] ? DMemory_697 : _GEN_789; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_791 = 10'h2ba == EXMEMALUOut[9:0] ? DMemory_698 : _GEN_790; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_792 = 10'h2bb == EXMEMALUOut[9:0] ? DMemory_699 : _GEN_791; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_793 = 10'h2bc == EXMEMALUOut[9:0] ? DMemory_700 : _GEN_792; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_794 = 10'h2bd == EXMEMALUOut[9:0] ? DMemory_701 : _GEN_793; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_795 = 10'h2be == EXMEMALUOut[9:0] ? DMemory_702 : _GEN_794; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_796 = 10'h2bf == EXMEMALUOut[9:0] ? DMemory_703 : _GEN_795; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_797 = 10'h2c0 == EXMEMALUOut[9:0] ? DMemory_704 : _GEN_796; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_798 = 10'h2c1 == EXMEMALUOut[9:0] ? DMemory_705 : _GEN_797; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_799 = 10'h2c2 == EXMEMALUOut[9:0] ? DMemory_706 : _GEN_798; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_800 = 10'h2c3 == EXMEMALUOut[9:0] ? DMemory_707 : _GEN_799; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_801 = 10'h2c4 == EXMEMALUOut[9:0] ? DMemory_708 : _GEN_800; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_802 = 10'h2c5 == EXMEMALUOut[9:0] ? DMemory_709 : _GEN_801; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_803 = 10'h2c6 == EXMEMALUOut[9:0] ? DMemory_710 : _GEN_802; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_804 = 10'h2c7 == EXMEMALUOut[9:0] ? DMemory_711 : _GEN_803; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_805 = 10'h2c8 == EXMEMALUOut[9:0] ? DMemory_712 : _GEN_804; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_806 = 10'h2c9 == EXMEMALUOut[9:0] ? DMemory_713 : _GEN_805; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_807 = 10'h2ca == EXMEMALUOut[9:0] ? DMemory_714 : _GEN_806; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_808 = 10'h2cb == EXMEMALUOut[9:0] ? DMemory_715 : _GEN_807; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_809 = 10'h2cc == EXMEMALUOut[9:0] ? DMemory_716 : _GEN_808; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_810 = 10'h2cd == EXMEMALUOut[9:0] ? DMemory_717 : _GEN_809; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_811 = 10'h2ce == EXMEMALUOut[9:0] ? DMemory_718 : _GEN_810; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_812 = 10'h2cf == EXMEMALUOut[9:0] ? DMemory_719 : _GEN_811; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_813 = 10'h2d0 == EXMEMALUOut[9:0] ? DMemory_720 : _GEN_812; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_814 = 10'h2d1 == EXMEMALUOut[9:0] ? DMemory_721 : _GEN_813; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_815 = 10'h2d2 == EXMEMALUOut[9:0] ? DMemory_722 : _GEN_814; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_816 = 10'h2d3 == EXMEMALUOut[9:0] ? DMemory_723 : _GEN_815; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_817 = 10'h2d4 == EXMEMALUOut[9:0] ? DMemory_724 : _GEN_816; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_818 = 10'h2d5 == EXMEMALUOut[9:0] ? DMemory_725 : _GEN_817; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_819 = 10'h2d6 == EXMEMALUOut[9:0] ? DMemory_726 : _GEN_818; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_820 = 10'h2d7 == EXMEMALUOut[9:0] ? DMemory_727 : _GEN_819; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_821 = 10'h2d8 == EXMEMALUOut[9:0] ? DMemory_728 : _GEN_820; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_822 = 10'h2d9 == EXMEMALUOut[9:0] ? DMemory_729 : _GEN_821; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_823 = 10'h2da == EXMEMALUOut[9:0] ? DMemory_730 : _GEN_822; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_824 = 10'h2db == EXMEMALUOut[9:0] ? DMemory_731 : _GEN_823; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_825 = 10'h2dc == EXMEMALUOut[9:0] ? DMemory_732 : _GEN_824; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_826 = 10'h2dd == EXMEMALUOut[9:0] ? DMemory_733 : _GEN_825; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_827 = 10'h2de == EXMEMALUOut[9:0] ? DMemory_734 : _GEN_826; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_828 = 10'h2df == EXMEMALUOut[9:0] ? DMemory_735 : _GEN_827; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_829 = 10'h2e0 == EXMEMALUOut[9:0] ? DMemory_736 : _GEN_828; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_830 = 10'h2e1 == EXMEMALUOut[9:0] ? DMemory_737 : _GEN_829; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_831 = 10'h2e2 == EXMEMALUOut[9:0] ? DMemory_738 : _GEN_830; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_832 = 10'h2e3 == EXMEMALUOut[9:0] ? DMemory_739 : _GEN_831; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_833 = 10'h2e4 == EXMEMALUOut[9:0] ? DMemory_740 : _GEN_832; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_834 = 10'h2e5 == EXMEMALUOut[9:0] ? DMemory_741 : _GEN_833; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_835 = 10'h2e6 == EXMEMALUOut[9:0] ? DMemory_742 : _GEN_834; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_836 = 10'h2e7 == EXMEMALUOut[9:0] ? DMemory_743 : _GEN_835; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_837 = 10'h2e8 == EXMEMALUOut[9:0] ? DMemory_744 : _GEN_836; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_838 = 10'h2e9 == EXMEMALUOut[9:0] ? DMemory_745 : _GEN_837; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_839 = 10'h2ea == EXMEMALUOut[9:0] ? DMemory_746 : _GEN_838; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_840 = 10'h2eb == EXMEMALUOut[9:0] ? DMemory_747 : _GEN_839; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_841 = 10'h2ec == EXMEMALUOut[9:0] ? DMemory_748 : _GEN_840; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_842 = 10'h2ed == EXMEMALUOut[9:0] ? DMemory_749 : _GEN_841; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_843 = 10'h2ee == EXMEMALUOut[9:0] ? DMemory_750 : _GEN_842; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_844 = 10'h2ef == EXMEMALUOut[9:0] ? DMemory_751 : _GEN_843; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_845 = 10'h2f0 == EXMEMALUOut[9:0] ? DMemory_752 : _GEN_844; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_846 = 10'h2f1 == EXMEMALUOut[9:0] ? DMemory_753 : _GEN_845; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_847 = 10'h2f2 == EXMEMALUOut[9:0] ? DMemory_754 : _GEN_846; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_848 = 10'h2f3 == EXMEMALUOut[9:0] ? DMemory_755 : _GEN_847; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_849 = 10'h2f4 == EXMEMALUOut[9:0] ? DMemory_756 : _GEN_848; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_850 = 10'h2f5 == EXMEMALUOut[9:0] ? DMemory_757 : _GEN_849; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_851 = 10'h2f6 == EXMEMALUOut[9:0] ? DMemory_758 : _GEN_850; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_852 = 10'h2f7 == EXMEMALUOut[9:0] ? DMemory_759 : _GEN_851; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_853 = 10'h2f8 == EXMEMALUOut[9:0] ? DMemory_760 : _GEN_852; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_854 = 10'h2f9 == EXMEMALUOut[9:0] ? DMemory_761 : _GEN_853; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_855 = 10'h2fa == EXMEMALUOut[9:0] ? DMemory_762 : _GEN_854; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_856 = 10'h2fb == EXMEMALUOut[9:0] ? DMemory_763 : _GEN_855; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_857 = 10'h2fc == EXMEMALUOut[9:0] ? DMemory_764 : _GEN_856; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_858 = 10'h2fd == EXMEMALUOut[9:0] ? DMemory_765 : _GEN_857; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_859 = 10'h2fe == EXMEMALUOut[9:0] ? DMemory_766 : _GEN_858; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_860 = 10'h2ff == EXMEMALUOut[9:0] ? DMemory_767 : _GEN_859; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_861 = 10'h300 == EXMEMALUOut[9:0] ? DMemory_768 : _GEN_860; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_862 = 10'h301 == EXMEMALUOut[9:0] ? DMemory_769 : _GEN_861; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_863 = 10'h302 == EXMEMALUOut[9:0] ? DMemory_770 : _GEN_862; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_864 = 10'h303 == EXMEMALUOut[9:0] ? DMemory_771 : _GEN_863; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_865 = 10'h304 == EXMEMALUOut[9:0] ? DMemory_772 : _GEN_864; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_866 = 10'h305 == EXMEMALUOut[9:0] ? DMemory_773 : _GEN_865; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_867 = 10'h306 == EXMEMALUOut[9:0] ? DMemory_774 : _GEN_866; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_868 = 10'h307 == EXMEMALUOut[9:0] ? DMemory_775 : _GEN_867; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_869 = 10'h308 == EXMEMALUOut[9:0] ? DMemory_776 : _GEN_868; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_870 = 10'h309 == EXMEMALUOut[9:0] ? DMemory_777 : _GEN_869; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_871 = 10'h30a == EXMEMALUOut[9:0] ? DMemory_778 : _GEN_870; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_872 = 10'h30b == EXMEMALUOut[9:0] ? DMemory_779 : _GEN_871; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_873 = 10'h30c == EXMEMALUOut[9:0] ? DMemory_780 : _GEN_872; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_874 = 10'h30d == EXMEMALUOut[9:0] ? DMemory_781 : _GEN_873; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_875 = 10'h30e == EXMEMALUOut[9:0] ? DMemory_782 : _GEN_874; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_876 = 10'h30f == EXMEMALUOut[9:0] ? DMemory_783 : _GEN_875; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_877 = 10'h310 == EXMEMALUOut[9:0] ? DMemory_784 : _GEN_876; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_878 = 10'h311 == EXMEMALUOut[9:0] ? DMemory_785 : _GEN_877; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_879 = 10'h312 == EXMEMALUOut[9:0] ? DMemory_786 : _GEN_878; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_880 = 10'h313 == EXMEMALUOut[9:0] ? DMemory_787 : _GEN_879; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_881 = 10'h314 == EXMEMALUOut[9:0] ? DMemory_788 : _GEN_880; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_882 = 10'h315 == EXMEMALUOut[9:0] ? DMemory_789 : _GEN_881; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_883 = 10'h316 == EXMEMALUOut[9:0] ? DMemory_790 : _GEN_882; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_884 = 10'h317 == EXMEMALUOut[9:0] ? DMemory_791 : _GEN_883; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_885 = 10'h318 == EXMEMALUOut[9:0] ? DMemory_792 : _GEN_884; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_886 = 10'h319 == EXMEMALUOut[9:0] ? DMemory_793 : _GEN_885; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_887 = 10'h31a == EXMEMALUOut[9:0] ? DMemory_794 : _GEN_886; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_888 = 10'h31b == EXMEMALUOut[9:0] ? DMemory_795 : _GEN_887; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_889 = 10'h31c == EXMEMALUOut[9:0] ? DMemory_796 : _GEN_888; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_890 = 10'h31d == EXMEMALUOut[9:0] ? DMemory_797 : _GEN_889; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_891 = 10'h31e == EXMEMALUOut[9:0] ? DMemory_798 : _GEN_890; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_892 = 10'h31f == EXMEMALUOut[9:0] ? DMemory_799 : _GEN_891; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_893 = 10'h320 == EXMEMALUOut[9:0] ? DMemory_800 : _GEN_892; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_894 = 10'h321 == EXMEMALUOut[9:0] ? DMemory_801 : _GEN_893; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_895 = 10'h322 == EXMEMALUOut[9:0] ? DMemory_802 : _GEN_894; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_896 = 10'h323 == EXMEMALUOut[9:0] ? DMemory_803 : _GEN_895; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_897 = 10'h324 == EXMEMALUOut[9:0] ? DMemory_804 : _GEN_896; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_898 = 10'h325 == EXMEMALUOut[9:0] ? DMemory_805 : _GEN_897; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_899 = 10'h326 == EXMEMALUOut[9:0] ? DMemory_806 : _GEN_898; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_900 = 10'h327 == EXMEMALUOut[9:0] ? DMemory_807 : _GEN_899; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_901 = 10'h328 == EXMEMALUOut[9:0] ? DMemory_808 : _GEN_900; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_902 = 10'h329 == EXMEMALUOut[9:0] ? DMemory_809 : _GEN_901; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_903 = 10'h32a == EXMEMALUOut[9:0] ? DMemory_810 : _GEN_902; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_904 = 10'h32b == EXMEMALUOut[9:0] ? DMemory_811 : _GEN_903; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_905 = 10'h32c == EXMEMALUOut[9:0] ? DMemory_812 : _GEN_904; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_906 = 10'h32d == EXMEMALUOut[9:0] ? DMemory_813 : _GEN_905; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_907 = 10'h32e == EXMEMALUOut[9:0] ? DMemory_814 : _GEN_906; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_908 = 10'h32f == EXMEMALUOut[9:0] ? DMemory_815 : _GEN_907; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_909 = 10'h330 == EXMEMALUOut[9:0] ? DMemory_816 : _GEN_908; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_910 = 10'h331 == EXMEMALUOut[9:0] ? DMemory_817 : _GEN_909; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_911 = 10'h332 == EXMEMALUOut[9:0] ? DMemory_818 : _GEN_910; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_912 = 10'h333 == EXMEMALUOut[9:0] ? DMemory_819 : _GEN_911; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_913 = 10'h334 == EXMEMALUOut[9:0] ? DMemory_820 : _GEN_912; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_914 = 10'h335 == EXMEMALUOut[9:0] ? DMemory_821 : _GEN_913; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_915 = 10'h336 == EXMEMALUOut[9:0] ? DMemory_822 : _GEN_914; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_916 = 10'h337 == EXMEMALUOut[9:0] ? DMemory_823 : _GEN_915; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_917 = 10'h338 == EXMEMALUOut[9:0] ? DMemory_824 : _GEN_916; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_918 = 10'h339 == EXMEMALUOut[9:0] ? DMemory_825 : _GEN_917; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_919 = 10'h33a == EXMEMALUOut[9:0] ? DMemory_826 : _GEN_918; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_920 = 10'h33b == EXMEMALUOut[9:0] ? DMemory_827 : _GEN_919; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_921 = 10'h33c == EXMEMALUOut[9:0] ? DMemory_828 : _GEN_920; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_922 = 10'h33d == EXMEMALUOut[9:0] ? DMemory_829 : _GEN_921; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_923 = 10'h33e == EXMEMALUOut[9:0] ? DMemory_830 : _GEN_922; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_924 = 10'h33f == EXMEMALUOut[9:0] ? DMemory_831 : _GEN_923; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_925 = 10'h340 == EXMEMALUOut[9:0] ? DMemory_832 : _GEN_924; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_926 = 10'h341 == EXMEMALUOut[9:0] ? DMemory_833 : _GEN_925; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_927 = 10'h342 == EXMEMALUOut[9:0] ? DMemory_834 : _GEN_926; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_928 = 10'h343 == EXMEMALUOut[9:0] ? DMemory_835 : _GEN_927; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_929 = 10'h344 == EXMEMALUOut[9:0] ? DMemory_836 : _GEN_928; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_930 = 10'h345 == EXMEMALUOut[9:0] ? DMemory_837 : _GEN_929; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_931 = 10'h346 == EXMEMALUOut[9:0] ? DMemory_838 : _GEN_930; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_932 = 10'h347 == EXMEMALUOut[9:0] ? DMemory_839 : _GEN_931; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_933 = 10'h348 == EXMEMALUOut[9:0] ? DMemory_840 : _GEN_932; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_934 = 10'h349 == EXMEMALUOut[9:0] ? DMemory_841 : _GEN_933; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_935 = 10'h34a == EXMEMALUOut[9:0] ? DMemory_842 : _GEN_934; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_936 = 10'h34b == EXMEMALUOut[9:0] ? DMemory_843 : _GEN_935; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_937 = 10'h34c == EXMEMALUOut[9:0] ? DMemory_844 : _GEN_936; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_938 = 10'h34d == EXMEMALUOut[9:0] ? DMemory_845 : _GEN_937; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_939 = 10'h34e == EXMEMALUOut[9:0] ? DMemory_846 : _GEN_938; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_940 = 10'h34f == EXMEMALUOut[9:0] ? DMemory_847 : _GEN_939; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_941 = 10'h350 == EXMEMALUOut[9:0] ? DMemory_848 : _GEN_940; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_942 = 10'h351 == EXMEMALUOut[9:0] ? DMemory_849 : _GEN_941; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_943 = 10'h352 == EXMEMALUOut[9:0] ? DMemory_850 : _GEN_942; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_944 = 10'h353 == EXMEMALUOut[9:0] ? DMemory_851 : _GEN_943; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_945 = 10'h354 == EXMEMALUOut[9:0] ? DMemory_852 : _GEN_944; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_946 = 10'h355 == EXMEMALUOut[9:0] ? DMemory_853 : _GEN_945; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_947 = 10'h356 == EXMEMALUOut[9:0] ? DMemory_854 : _GEN_946; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_948 = 10'h357 == EXMEMALUOut[9:0] ? DMemory_855 : _GEN_947; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_949 = 10'h358 == EXMEMALUOut[9:0] ? DMemory_856 : _GEN_948; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_950 = 10'h359 == EXMEMALUOut[9:0] ? DMemory_857 : _GEN_949; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_951 = 10'h35a == EXMEMALUOut[9:0] ? DMemory_858 : _GEN_950; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_952 = 10'h35b == EXMEMALUOut[9:0] ? DMemory_859 : _GEN_951; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_953 = 10'h35c == EXMEMALUOut[9:0] ? DMemory_860 : _GEN_952; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_954 = 10'h35d == EXMEMALUOut[9:0] ? DMemory_861 : _GEN_953; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_955 = 10'h35e == EXMEMALUOut[9:0] ? DMemory_862 : _GEN_954; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_956 = 10'h35f == EXMEMALUOut[9:0] ? DMemory_863 : _GEN_955; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_957 = 10'h360 == EXMEMALUOut[9:0] ? DMemory_864 : _GEN_956; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_958 = 10'h361 == EXMEMALUOut[9:0] ? DMemory_865 : _GEN_957; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_959 = 10'h362 == EXMEMALUOut[9:0] ? DMemory_866 : _GEN_958; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_960 = 10'h363 == EXMEMALUOut[9:0] ? DMemory_867 : _GEN_959; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_961 = 10'h364 == EXMEMALUOut[9:0] ? DMemory_868 : _GEN_960; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_962 = 10'h365 == EXMEMALUOut[9:0] ? DMemory_869 : _GEN_961; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_963 = 10'h366 == EXMEMALUOut[9:0] ? DMemory_870 : _GEN_962; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_964 = 10'h367 == EXMEMALUOut[9:0] ? DMemory_871 : _GEN_963; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_965 = 10'h368 == EXMEMALUOut[9:0] ? DMemory_872 : _GEN_964; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_966 = 10'h369 == EXMEMALUOut[9:0] ? DMemory_873 : _GEN_965; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_967 = 10'h36a == EXMEMALUOut[9:0] ? DMemory_874 : _GEN_966; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_968 = 10'h36b == EXMEMALUOut[9:0] ? DMemory_875 : _GEN_967; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_969 = 10'h36c == EXMEMALUOut[9:0] ? DMemory_876 : _GEN_968; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_970 = 10'h36d == EXMEMALUOut[9:0] ? DMemory_877 : _GEN_969; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_971 = 10'h36e == EXMEMALUOut[9:0] ? DMemory_878 : _GEN_970; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_972 = 10'h36f == EXMEMALUOut[9:0] ? DMemory_879 : _GEN_971; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_973 = 10'h370 == EXMEMALUOut[9:0] ? DMemory_880 : _GEN_972; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_974 = 10'h371 == EXMEMALUOut[9:0] ? DMemory_881 : _GEN_973; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_975 = 10'h372 == EXMEMALUOut[9:0] ? DMemory_882 : _GEN_974; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_976 = 10'h373 == EXMEMALUOut[9:0] ? DMemory_883 : _GEN_975; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_977 = 10'h374 == EXMEMALUOut[9:0] ? DMemory_884 : _GEN_976; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_978 = 10'h375 == EXMEMALUOut[9:0] ? DMemory_885 : _GEN_977; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_979 = 10'h376 == EXMEMALUOut[9:0] ? DMemory_886 : _GEN_978; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_980 = 10'h377 == EXMEMALUOut[9:0] ? DMemory_887 : _GEN_979; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_981 = 10'h378 == EXMEMALUOut[9:0] ? DMemory_888 : _GEN_980; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_982 = 10'h379 == EXMEMALUOut[9:0] ? DMemory_889 : _GEN_981; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_983 = 10'h37a == EXMEMALUOut[9:0] ? DMemory_890 : _GEN_982; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_984 = 10'h37b == EXMEMALUOut[9:0] ? DMemory_891 : _GEN_983; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_985 = 10'h37c == EXMEMALUOut[9:0] ? DMemory_892 : _GEN_984; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_986 = 10'h37d == EXMEMALUOut[9:0] ? DMemory_893 : _GEN_985; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_987 = 10'h37e == EXMEMALUOut[9:0] ? DMemory_894 : _GEN_986; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_988 = 10'h37f == EXMEMALUOut[9:0] ? DMemory_895 : _GEN_987; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_989 = 10'h380 == EXMEMALUOut[9:0] ? DMemory_896 : _GEN_988; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_990 = 10'h381 == EXMEMALUOut[9:0] ? DMemory_897 : _GEN_989; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_991 = 10'h382 == EXMEMALUOut[9:0] ? DMemory_898 : _GEN_990; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_992 = 10'h383 == EXMEMALUOut[9:0] ? DMemory_899 : _GEN_991; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_993 = 10'h384 == EXMEMALUOut[9:0] ? DMemory_900 : _GEN_992; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_994 = 10'h385 == EXMEMALUOut[9:0] ? DMemory_901 : _GEN_993; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_995 = 10'h386 == EXMEMALUOut[9:0] ? DMemory_902 : _GEN_994; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_996 = 10'h387 == EXMEMALUOut[9:0] ? DMemory_903 : _GEN_995; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_997 = 10'h388 == EXMEMALUOut[9:0] ? DMemory_904 : _GEN_996; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_998 = 10'h389 == EXMEMALUOut[9:0] ? DMemory_905 : _GEN_997; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_999 = 10'h38a == EXMEMALUOut[9:0] ? DMemory_906 : _GEN_998; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1000 = 10'h38b == EXMEMALUOut[9:0] ? DMemory_907 : _GEN_999; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1001 = 10'h38c == EXMEMALUOut[9:0] ? DMemory_908 : _GEN_1000; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1002 = 10'h38d == EXMEMALUOut[9:0] ? DMemory_909 : _GEN_1001; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1003 = 10'h38e == EXMEMALUOut[9:0] ? DMemory_910 : _GEN_1002; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1004 = 10'h38f == EXMEMALUOut[9:0] ? DMemory_911 : _GEN_1003; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1005 = 10'h390 == EXMEMALUOut[9:0] ? DMemory_912 : _GEN_1004; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1006 = 10'h391 == EXMEMALUOut[9:0] ? DMemory_913 : _GEN_1005; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1007 = 10'h392 == EXMEMALUOut[9:0] ? DMemory_914 : _GEN_1006; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1008 = 10'h393 == EXMEMALUOut[9:0] ? DMemory_915 : _GEN_1007; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1009 = 10'h394 == EXMEMALUOut[9:0] ? DMemory_916 : _GEN_1008; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1010 = 10'h395 == EXMEMALUOut[9:0] ? DMemory_917 : _GEN_1009; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1011 = 10'h396 == EXMEMALUOut[9:0] ? DMemory_918 : _GEN_1010; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1012 = 10'h397 == EXMEMALUOut[9:0] ? DMemory_919 : _GEN_1011; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1013 = 10'h398 == EXMEMALUOut[9:0] ? DMemory_920 : _GEN_1012; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1014 = 10'h399 == EXMEMALUOut[9:0] ? DMemory_921 : _GEN_1013; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1015 = 10'h39a == EXMEMALUOut[9:0] ? DMemory_922 : _GEN_1014; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1016 = 10'h39b == EXMEMALUOut[9:0] ? DMemory_923 : _GEN_1015; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1017 = 10'h39c == EXMEMALUOut[9:0] ? DMemory_924 : _GEN_1016; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1018 = 10'h39d == EXMEMALUOut[9:0] ? DMemory_925 : _GEN_1017; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1019 = 10'h39e == EXMEMALUOut[9:0] ? DMemory_926 : _GEN_1018; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1020 = 10'h39f == EXMEMALUOut[9:0] ? DMemory_927 : _GEN_1019; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1021 = 10'h3a0 == EXMEMALUOut[9:0] ? DMemory_928 : _GEN_1020; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1022 = 10'h3a1 == EXMEMALUOut[9:0] ? DMemory_929 : _GEN_1021; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1023 = 10'h3a2 == EXMEMALUOut[9:0] ? DMemory_930 : _GEN_1022; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1024 = 10'h3a3 == EXMEMALUOut[9:0] ? DMemory_931 : _GEN_1023; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1025 = 10'h3a4 == EXMEMALUOut[9:0] ? DMemory_932 : _GEN_1024; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1026 = 10'h3a5 == EXMEMALUOut[9:0] ? DMemory_933 : _GEN_1025; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1027 = 10'h3a6 == EXMEMALUOut[9:0] ? DMemory_934 : _GEN_1026; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1028 = 10'h3a7 == EXMEMALUOut[9:0] ? DMemory_935 : _GEN_1027; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1029 = 10'h3a8 == EXMEMALUOut[9:0] ? DMemory_936 : _GEN_1028; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1030 = 10'h3a9 == EXMEMALUOut[9:0] ? DMemory_937 : _GEN_1029; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1031 = 10'h3aa == EXMEMALUOut[9:0] ? DMemory_938 : _GEN_1030; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1032 = 10'h3ab == EXMEMALUOut[9:0] ? DMemory_939 : _GEN_1031; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1033 = 10'h3ac == EXMEMALUOut[9:0] ? DMemory_940 : _GEN_1032; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1034 = 10'h3ad == EXMEMALUOut[9:0] ? DMemory_941 : _GEN_1033; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1035 = 10'h3ae == EXMEMALUOut[9:0] ? DMemory_942 : _GEN_1034; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1036 = 10'h3af == EXMEMALUOut[9:0] ? DMemory_943 : _GEN_1035; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1037 = 10'h3b0 == EXMEMALUOut[9:0] ? DMemory_944 : _GEN_1036; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1038 = 10'h3b1 == EXMEMALUOut[9:0] ? DMemory_945 : _GEN_1037; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1039 = 10'h3b2 == EXMEMALUOut[9:0] ? DMemory_946 : _GEN_1038; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1040 = 10'h3b3 == EXMEMALUOut[9:0] ? DMemory_947 : _GEN_1039; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1041 = 10'h3b4 == EXMEMALUOut[9:0] ? DMemory_948 : _GEN_1040; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1042 = 10'h3b5 == EXMEMALUOut[9:0] ? DMemory_949 : _GEN_1041; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1043 = 10'h3b6 == EXMEMALUOut[9:0] ? DMemory_950 : _GEN_1042; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1044 = 10'h3b7 == EXMEMALUOut[9:0] ? DMemory_951 : _GEN_1043; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1045 = 10'h3b8 == EXMEMALUOut[9:0] ? DMemory_952 : _GEN_1044; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1046 = 10'h3b9 == EXMEMALUOut[9:0] ? DMemory_953 : _GEN_1045; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1047 = 10'h3ba == EXMEMALUOut[9:0] ? DMemory_954 : _GEN_1046; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1048 = 10'h3bb == EXMEMALUOut[9:0] ? DMemory_955 : _GEN_1047; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1049 = 10'h3bc == EXMEMALUOut[9:0] ? DMemory_956 : _GEN_1048; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1050 = 10'h3bd == EXMEMALUOut[9:0] ? DMemory_957 : _GEN_1049; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1051 = 10'h3be == EXMEMALUOut[9:0] ? DMemory_958 : _GEN_1050; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1052 = 10'h3bf == EXMEMALUOut[9:0] ? DMemory_959 : _GEN_1051; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1053 = 10'h3c0 == EXMEMALUOut[9:0] ? DMemory_960 : _GEN_1052; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1054 = 10'h3c1 == EXMEMALUOut[9:0] ? DMemory_961 : _GEN_1053; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1055 = 10'h3c2 == EXMEMALUOut[9:0] ? DMemory_962 : _GEN_1054; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1056 = 10'h3c3 == EXMEMALUOut[9:0] ? DMemory_963 : _GEN_1055; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1057 = 10'h3c4 == EXMEMALUOut[9:0] ? DMemory_964 : _GEN_1056; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1058 = 10'h3c5 == EXMEMALUOut[9:0] ? DMemory_965 : _GEN_1057; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1059 = 10'h3c6 == EXMEMALUOut[9:0] ? DMemory_966 : _GEN_1058; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1060 = 10'h3c7 == EXMEMALUOut[9:0] ? DMemory_967 : _GEN_1059; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1061 = 10'h3c8 == EXMEMALUOut[9:0] ? DMemory_968 : _GEN_1060; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1062 = 10'h3c9 == EXMEMALUOut[9:0] ? DMemory_969 : _GEN_1061; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1063 = 10'h3ca == EXMEMALUOut[9:0] ? DMemory_970 : _GEN_1062; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1064 = 10'h3cb == EXMEMALUOut[9:0] ? DMemory_971 : _GEN_1063; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1065 = 10'h3cc == EXMEMALUOut[9:0] ? DMemory_972 : _GEN_1064; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1066 = 10'h3cd == EXMEMALUOut[9:0] ? DMemory_973 : _GEN_1065; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1067 = 10'h3ce == EXMEMALUOut[9:0] ? DMemory_974 : _GEN_1066; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1068 = 10'h3cf == EXMEMALUOut[9:0] ? DMemory_975 : _GEN_1067; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1069 = 10'h3d0 == EXMEMALUOut[9:0] ? DMemory_976 : _GEN_1068; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1070 = 10'h3d1 == EXMEMALUOut[9:0] ? DMemory_977 : _GEN_1069; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1071 = 10'h3d2 == EXMEMALUOut[9:0] ? DMemory_978 : _GEN_1070; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1072 = 10'h3d3 == EXMEMALUOut[9:0] ? DMemory_979 : _GEN_1071; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1073 = 10'h3d4 == EXMEMALUOut[9:0] ? DMemory_980 : _GEN_1072; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1074 = 10'h3d5 == EXMEMALUOut[9:0] ? DMemory_981 : _GEN_1073; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1075 = 10'h3d6 == EXMEMALUOut[9:0] ? DMemory_982 : _GEN_1074; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1076 = 10'h3d7 == EXMEMALUOut[9:0] ? DMemory_983 : _GEN_1075; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1077 = 10'h3d8 == EXMEMALUOut[9:0] ? DMemory_984 : _GEN_1076; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1078 = 10'h3d9 == EXMEMALUOut[9:0] ? DMemory_985 : _GEN_1077; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1079 = 10'h3da == EXMEMALUOut[9:0] ? DMemory_986 : _GEN_1078; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1080 = 10'h3db == EXMEMALUOut[9:0] ? DMemory_987 : _GEN_1079; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1081 = 10'h3dc == EXMEMALUOut[9:0] ? DMemory_988 : _GEN_1080; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1082 = 10'h3dd == EXMEMALUOut[9:0] ? DMemory_989 : _GEN_1081; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1083 = 10'h3de == EXMEMALUOut[9:0] ? DMemory_990 : _GEN_1082; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1084 = 10'h3df == EXMEMALUOut[9:0] ? DMemory_991 : _GEN_1083; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1085 = 10'h3e0 == EXMEMALUOut[9:0] ? DMemory_992 : _GEN_1084; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1086 = 10'h3e1 == EXMEMALUOut[9:0] ? DMemory_993 : _GEN_1085; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1087 = 10'h3e2 == EXMEMALUOut[9:0] ? DMemory_994 : _GEN_1086; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1088 = 10'h3e3 == EXMEMALUOut[9:0] ? DMemory_995 : _GEN_1087; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1089 = 10'h3e4 == EXMEMALUOut[9:0] ? DMemory_996 : _GEN_1088; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1090 = 10'h3e5 == EXMEMALUOut[9:0] ? DMemory_997 : _GEN_1089; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1091 = 10'h3e6 == EXMEMALUOut[9:0] ? DMemory_998 : _GEN_1090; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1092 = 10'h3e7 == EXMEMALUOut[9:0] ? DMemory_999 : _GEN_1091; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1093 = 10'h3e8 == EXMEMALUOut[9:0] ? DMemory_1000 : _GEN_1092; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1094 = 10'h3e9 == EXMEMALUOut[9:0] ? DMemory_1001 : _GEN_1093; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1095 = 10'h3ea == EXMEMALUOut[9:0] ? DMemory_1002 : _GEN_1094; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1096 = 10'h3eb == EXMEMALUOut[9:0] ? DMemory_1003 : _GEN_1095; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1097 = 10'h3ec == EXMEMALUOut[9:0] ? DMemory_1004 : _GEN_1096; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1098 = 10'h3ed == EXMEMALUOut[9:0] ? DMemory_1005 : _GEN_1097; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1099 = 10'h3ee == EXMEMALUOut[9:0] ? DMemory_1006 : _GEN_1098; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1100 = 10'h3ef == EXMEMALUOut[9:0] ? DMemory_1007 : _GEN_1099; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1101 = 10'h3f0 == EXMEMALUOut[9:0] ? DMemory_1008 : _GEN_1100; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1102 = 10'h3f1 == EXMEMALUOut[9:0] ? DMemory_1009 : _GEN_1101; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1103 = 10'h3f2 == EXMEMALUOut[9:0] ? DMemory_1010 : _GEN_1102; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1104 = 10'h3f3 == EXMEMALUOut[9:0] ? DMemory_1011 : _GEN_1103; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1105 = 10'h3f4 == EXMEMALUOut[9:0] ? DMemory_1012 : _GEN_1104; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1106 = 10'h3f5 == EXMEMALUOut[9:0] ? DMemory_1013 : _GEN_1105; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1107 = 10'h3f6 == EXMEMALUOut[9:0] ? DMemory_1014 : _GEN_1106; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1108 = 10'h3f7 == EXMEMALUOut[9:0] ? DMemory_1015 : _GEN_1107; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1109 = 10'h3f8 == EXMEMALUOut[9:0] ? DMemory_1016 : _GEN_1108; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1110 = 10'h3f9 == EXMEMALUOut[9:0] ? DMemory_1017 : _GEN_1109; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1111 = 10'h3fa == EXMEMALUOut[9:0] ? DMemory_1018 : _GEN_1110; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1112 = 10'h3fb == EXMEMALUOut[9:0] ? DMemory_1019 : _GEN_1111; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1113 = 10'h3fc == EXMEMALUOut[9:0] ? DMemory_1020 : _GEN_1112; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1114 = 10'h3fd == EXMEMALUOut[9:0] ? DMemory_1021 : _GEN_1113; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1115 = 10'h3fe == EXMEMALUOut[9:0] ? DMemory_1022 : _GEN_1114; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1116 = 10'h3ff == EXMEMALUOut[9:0] ? DMemory_1023 : _GEN_1115; // @[cpu.scala 435:{18,18}]
  wire [31:0] _GEN_1117 = 10'h0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_0; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1118 = 10'h1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1119 = 10'h2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_2; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1120 = 10'h3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_3; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1121 = 10'h4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_4; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1122 = 10'h5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_5; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1123 = 10'h6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_6; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1124 = 10'h7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_7; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1125 = 10'h8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_8; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1126 = 10'h9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_9; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1127 = 10'ha == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_10; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1128 = 10'hb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_11; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1129 = 10'hc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_12; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1130 = 10'hd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_13; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1131 = 10'he == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_14; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1132 = 10'hf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_15; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1133 = 10'h10 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_16; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1134 = 10'h11 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_17; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1135 = 10'h12 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_18; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1136 = 10'h13 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_19; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1137 = 10'h14 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_20; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1138 = 10'h15 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_21; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1139 = 10'h16 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_22; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1140 = 10'h17 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_23; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1141 = 10'h18 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_24; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1142 = 10'h19 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_25; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1143 = 10'h1a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_26; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1144 = 10'h1b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_27; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1145 = 10'h1c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_28; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1146 = 10'h1d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_29; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1147 = 10'h1e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_30; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1148 = 10'h1f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_31; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1149 = 10'h20 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_32; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1150 = 10'h21 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_33; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1151 = 10'h22 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_34; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1152 = 10'h23 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_35; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1153 = 10'h24 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_36; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1154 = 10'h25 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_37; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1155 = 10'h26 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_38; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1156 = 10'h27 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_39; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1157 = 10'h28 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_40; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1158 = 10'h29 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_41; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1159 = 10'h2a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_42; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1160 = 10'h2b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_43; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1161 = 10'h2c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_44; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1162 = 10'h2d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_45; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1163 = 10'h2e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_46; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1164 = 10'h2f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_47; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1165 = 10'h30 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_48; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1166 = 10'h31 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_49; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1167 = 10'h32 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_50; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1168 = 10'h33 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_51; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1169 = 10'h34 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_52; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1170 = 10'h35 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_53; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1171 = 10'h36 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_54; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1172 = 10'h37 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_55; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1173 = 10'h38 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_56; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1174 = 10'h39 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_57; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1175 = 10'h3a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_58; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1176 = 10'h3b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_59; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1177 = 10'h3c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_60; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1178 = 10'h3d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_61; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1179 = 10'h3e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_62; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1180 = 10'h3f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_63; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1181 = 10'h40 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_64; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1182 = 10'h41 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_65; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1183 = 10'h42 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_66; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1184 = 10'h43 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_67; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1185 = 10'h44 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_68; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1186 = 10'h45 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_69; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1187 = 10'h46 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_70; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1188 = 10'h47 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_71; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1189 = 10'h48 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_72; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1190 = 10'h49 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_73; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1191 = 10'h4a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_74; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1192 = 10'h4b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_75; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1193 = 10'h4c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_76; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1194 = 10'h4d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_77; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1195 = 10'h4e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_78; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1196 = 10'h4f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_79; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1197 = 10'h50 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_80; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1198 = 10'h51 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_81; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1199 = 10'h52 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_82; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1200 = 10'h53 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_83; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1201 = 10'h54 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_84; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1202 = 10'h55 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_85; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1203 = 10'h56 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_86; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1204 = 10'h57 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_87; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1205 = 10'h58 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_88; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1206 = 10'h59 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_89; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1207 = 10'h5a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_90; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1208 = 10'h5b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_91; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1209 = 10'h5c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_92; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1210 = 10'h5d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_93; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1211 = 10'h5e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_94; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1212 = 10'h5f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_95; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1213 = 10'h60 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_96; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1214 = 10'h61 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_97; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1215 = 10'h62 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_98; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1216 = 10'h63 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_99; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1217 = 10'h64 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_100; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1218 = 10'h65 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_101; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1219 = 10'h66 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_102; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1220 = 10'h67 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_103; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1221 = 10'h68 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_104; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1222 = 10'h69 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_105; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1223 = 10'h6a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_106; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1224 = 10'h6b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_107; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1225 = 10'h6c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_108; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1226 = 10'h6d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_109; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1227 = 10'h6e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_110; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1228 = 10'h6f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_111; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1229 = 10'h70 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_112; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1230 = 10'h71 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_113; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1231 = 10'h72 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_114; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1232 = 10'h73 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_115; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1233 = 10'h74 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_116; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1234 = 10'h75 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_117; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1235 = 10'h76 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_118; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1236 = 10'h77 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_119; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1237 = 10'h78 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_120; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1238 = 10'h79 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_121; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1239 = 10'h7a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_122; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1240 = 10'h7b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_123; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1241 = 10'h7c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_124; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1242 = 10'h7d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_125; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1243 = 10'h7e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_126; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1244 = 10'h7f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_127; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1245 = 10'h80 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_128; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1246 = 10'h81 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_129; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1247 = 10'h82 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_130; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1248 = 10'h83 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_131; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1249 = 10'h84 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_132; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1250 = 10'h85 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_133; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1251 = 10'h86 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_134; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1252 = 10'h87 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_135; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1253 = 10'h88 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_136; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1254 = 10'h89 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_137; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1255 = 10'h8a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_138; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1256 = 10'h8b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_139; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1257 = 10'h8c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_140; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1258 = 10'h8d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_141; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1259 = 10'h8e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_142; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1260 = 10'h8f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_143; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1261 = 10'h90 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_144; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1262 = 10'h91 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_145; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1263 = 10'h92 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_146; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1264 = 10'h93 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_147; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1265 = 10'h94 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_148; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1266 = 10'h95 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_149; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1267 = 10'h96 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_150; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1268 = 10'h97 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_151; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1269 = 10'h98 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_152; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1270 = 10'h99 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_153; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1271 = 10'h9a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_154; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1272 = 10'h9b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_155; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1273 = 10'h9c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_156; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1274 = 10'h9d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_157; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1275 = 10'h9e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_158; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1276 = 10'h9f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_159; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1277 = 10'ha0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_160; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1278 = 10'ha1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_161; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1279 = 10'ha2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_162; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1280 = 10'ha3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_163; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1281 = 10'ha4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_164; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1282 = 10'ha5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_165; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1283 = 10'ha6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_166; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1284 = 10'ha7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_167; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1285 = 10'ha8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_168; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1286 = 10'ha9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_169; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1287 = 10'haa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_170; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1288 = 10'hab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_171; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1289 = 10'hac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_172; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1290 = 10'had == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_173; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1291 = 10'hae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_174; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1292 = 10'haf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_175; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1293 = 10'hb0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_176; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1294 = 10'hb1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_177; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1295 = 10'hb2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_178; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1296 = 10'hb3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_179; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1297 = 10'hb4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_180; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1298 = 10'hb5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_181; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1299 = 10'hb6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_182; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1300 = 10'hb7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_183; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1301 = 10'hb8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_184; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1302 = 10'hb9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_185; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1303 = 10'hba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_186; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1304 = 10'hbb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_187; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1305 = 10'hbc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_188; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1306 = 10'hbd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_189; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1307 = 10'hbe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_190; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1308 = 10'hbf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_191; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1309 = 10'hc0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_192; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1310 = 10'hc1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_193; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1311 = 10'hc2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_194; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1312 = 10'hc3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_195; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1313 = 10'hc4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_196; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1314 = 10'hc5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_197; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1315 = 10'hc6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_198; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1316 = 10'hc7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_199; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1317 = 10'hc8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_200; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1318 = 10'hc9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_201; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1319 = 10'hca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_202; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1320 = 10'hcb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_203; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1321 = 10'hcc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_204; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1322 = 10'hcd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_205; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1323 = 10'hce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_206; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1324 = 10'hcf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_207; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1325 = 10'hd0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_208; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1326 = 10'hd1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_209; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1327 = 10'hd2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_210; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1328 = 10'hd3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_211; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1329 = 10'hd4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_212; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1330 = 10'hd5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_213; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1331 = 10'hd6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_214; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1332 = 10'hd7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_215; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1333 = 10'hd8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_216; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1334 = 10'hd9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_217; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1335 = 10'hda == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_218; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1336 = 10'hdb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_219; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1337 = 10'hdc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_220; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1338 = 10'hdd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_221; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1339 = 10'hde == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_222; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1340 = 10'hdf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_223; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1341 = 10'he0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_224; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1342 = 10'he1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_225; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1343 = 10'he2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_226; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1344 = 10'he3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_227; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1345 = 10'he4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_228; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1346 = 10'he5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_229; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1347 = 10'he6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_230; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1348 = 10'he7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_231; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1349 = 10'he8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_232; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1350 = 10'he9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_233; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1351 = 10'hea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_234; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1352 = 10'heb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_235; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1353 = 10'hec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_236; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1354 = 10'hed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_237; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1355 = 10'hee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_238; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1356 = 10'hef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_239; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1357 = 10'hf0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_240; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1358 = 10'hf1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_241; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1359 = 10'hf2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_242; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1360 = 10'hf3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_243; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1361 = 10'hf4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_244; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1362 = 10'hf5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_245; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1363 = 10'hf6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_246; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1364 = 10'hf7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_247; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1365 = 10'hf8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_248; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1366 = 10'hf9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_249; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1367 = 10'hfa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_250; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1368 = 10'hfb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_251; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1369 = 10'hfc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_252; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1370 = 10'hfd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_253; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1371 = 10'hfe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_254; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1372 = 10'hff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_255; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1373 = 10'h100 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_256; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1374 = 10'h101 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_257; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1375 = 10'h102 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_258; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1376 = 10'h103 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_259; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1377 = 10'h104 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_260; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1378 = 10'h105 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_261; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1379 = 10'h106 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_262; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1380 = 10'h107 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_263; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1381 = 10'h108 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_264; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1382 = 10'h109 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_265; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1383 = 10'h10a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_266; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1384 = 10'h10b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_267; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1385 = 10'h10c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_268; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1386 = 10'h10d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_269; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1387 = 10'h10e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_270; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1388 = 10'h10f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_271; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1389 = 10'h110 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_272; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1390 = 10'h111 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_273; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1391 = 10'h112 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_274; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1392 = 10'h113 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_275; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1393 = 10'h114 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_276; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1394 = 10'h115 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_277; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1395 = 10'h116 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_278; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1396 = 10'h117 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_279; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1397 = 10'h118 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_280; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1398 = 10'h119 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_281; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1399 = 10'h11a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_282; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1400 = 10'h11b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_283; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1401 = 10'h11c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_284; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1402 = 10'h11d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_285; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1403 = 10'h11e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_286; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1404 = 10'h11f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_287; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1405 = 10'h120 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_288; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1406 = 10'h121 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_289; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1407 = 10'h122 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_290; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1408 = 10'h123 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_291; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1409 = 10'h124 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_292; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1410 = 10'h125 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_293; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1411 = 10'h126 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_294; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1412 = 10'h127 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_295; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1413 = 10'h128 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_296; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1414 = 10'h129 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_297; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1415 = 10'h12a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_298; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1416 = 10'h12b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_299; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1417 = 10'h12c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_300; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1418 = 10'h12d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_301; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1419 = 10'h12e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_302; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1420 = 10'h12f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_303; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1421 = 10'h130 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_304; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1422 = 10'h131 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_305; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1423 = 10'h132 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_306; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1424 = 10'h133 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_307; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1425 = 10'h134 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_308; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1426 = 10'h135 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_309; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1427 = 10'h136 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_310; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1428 = 10'h137 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_311; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1429 = 10'h138 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_312; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1430 = 10'h139 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_313; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1431 = 10'h13a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_314; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1432 = 10'h13b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_315; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1433 = 10'h13c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_316; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1434 = 10'h13d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_317; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1435 = 10'h13e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_318; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1436 = 10'h13f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_319; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1437 = 10'h140 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_320; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1438 = 10'h141 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_321; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1439 = 10'h142 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_322; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1440 = 10'h143 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_323; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1441 = 10'h144 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_324; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1442 = 10'h145 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_325; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1443 = 10'h146 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_326; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1444 = 10'h147 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_327; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1445 = 10'h148 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_328; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1446 = 10'h149 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_329; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1447 = 10'h14a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_330; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1448 = 10'h14b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_331; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1449 = 10'h14c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_332; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1450 = 10'h14d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_333; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1451 = 10'h14e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_334; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1452 = 10'h14f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_335; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1453 = 10'h150 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_336; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1454 = 10'h151 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_337; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1455 = 10'h152 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_338; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1456 = 10'h153 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_339; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1457 = 10'h154 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_340; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1458 = 10'h155 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_341; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1459 = 10'h156 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_342; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1460 = 10'h157 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_343; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1461 = 10'h158 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_344; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1462 = 10'h159 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_345; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1463 = 10'h15a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_346; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1464 = 10'h15b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_347; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1465 = 10'h15c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_348; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1466 = 10'h15d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_349; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1467 = 10'h15e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_350; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1468 = 10'h15f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_351; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1469 = 10'h160 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_352; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1470 = 10'h161 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_353; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1471 = 10'h162 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_354; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1472 = 10'h163 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_355; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1473 = 10'h164 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_356; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1474 = 10'h165 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_357; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1475 = 10'h166 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_358; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1476 = 10'h167 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_359; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1477 = 10'h168 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_360; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1478 = 10'h169 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_361; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1479 = 10'h16a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_362; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1480 = 10'h16b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_363; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1481 = 10'h16c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_364; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1482 = 10'h16d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_365; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1483 = 10'h16e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_366; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1484 = 10'h16f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_367; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1485 = 10'h170 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_368; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1486 = 10'h171 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_369; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1487 = 10'h172 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_370; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1488 = 10'h173 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_371; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1489 = 10'h174 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_372; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1490 = 10'h175 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_373; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1491 = 10'h176 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_374; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1492 = 10'h177 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_375; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1493 = 10'h178 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_376; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1494 = 10'h179 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_377; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1495 = 10'h17a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_378; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1496 = 10'h17b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_379; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1497 = 10'h17c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_380; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1498 = 10'h17d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_381; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1499 = 10'h17e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_382; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1500 = 10'h17f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_383; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1501 = 10'h180 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_384; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1502 = 10'h181 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_385; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1503 = 10'h182 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_386; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1504 = 10'h183 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_387; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1505 = 10'h184 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_388; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1506 = 10'h185 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_389; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1507 = 10'h186 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_390; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1508 = 10'h187 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_391; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1509 = 10'h188 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_392; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1510 = 10'h189 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_393; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1511 = 10'h18a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_394; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1512 = 10'h18b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_395; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1513 = 10'h18c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_396; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1514 = 10'h18d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_397; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1515 = 10'h18e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_398; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1516 = 10'h18f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_399; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1517 = 10'h190 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_400; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1518 = 10'h191 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_401; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1519 = 10'h192 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_402; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1520 = 10'h193 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_403; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1521 = 10'h194 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_404; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1522 = 10'h195 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_405; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1523 = 10'h196 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_406; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1524 = 10'h197 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_407; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1525 = 10'h198 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_408; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1526 = 10'h199 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_409; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1527 = 10'h19a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_410; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1528 = 10'h19b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_411; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1529 = 10'h19c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_412; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1530 = 10'h19d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_413; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1531 = 10'h19e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_414; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1532 = 10'h19f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_415; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1533 = 10'h1a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_416; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1534 = 10'h1a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_417; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1535 = 10'h1a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_418; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1536 = 10'h1a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_419; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1537 = 10'h1a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_420; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1538 = 10'h1a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_421; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1539 = 10'h1a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_422; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1540 = 10'h1a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_423; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1541 = 10'h1a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_424; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1542 = 10'h1a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_425; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1543 = 10'h1aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_426; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1544 = 10'h1ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_427; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1545 = 10'h1ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_428; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1546 = 10'h1ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_429; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1547 = 10'h1ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_430; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1548 = 10'h1af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_431; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1549 = 10'h1b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_432; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1550 = 10'h1b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_433; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1551 = 10'h1b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_434; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1552 = 10'h1b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_435; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1553 = 10'h1b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_436; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1554 = 10'h1b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_437; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1555 = 10'h1b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_438; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1556 = 10'h1b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_439; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1557 = 10'h1b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_440; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1558 = 10'h1b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_441; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1559 = 10'h1ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_442; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1560 = 10'h1bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_443; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1561 = 10'h1bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_444; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1562 = 10'h1bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_445; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1563 = 10'h1be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_446; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1564 = 10'h1bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_447; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1565 = 10'h1c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_448; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1566 = 10'h1c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_449; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1567 = 10'h1c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_450; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1568 = 10'h1c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_451; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1569 = 10'h1c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_452; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1570 = 10'h1c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_453; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1571 = 10'h1c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_454; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1572 = 10'h1c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_455; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1573 = 10'h1c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_456; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1574 = 10'h1c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_457; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1575 = 10'h1ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_458; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1576 = 10'h1cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_459; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1577 = 10'h1cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_460; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1578 = 10'h1cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_461; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1579 = 10'h1ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_462; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1580 = 10'h1cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_463; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1581 = 10'h1d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_464; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1582 = 10'h1d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_465; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1583 = 10'h1d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_466; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1584 = 10'h1d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_467; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1585 = 10'h1d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_468; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1586 = 10'h1d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_469; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1587 = 10'h1d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_470; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1588 = 10'h1d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_471; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1589 = 10'h1d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_472; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1590 = 10'h1d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_473; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1591 = 10'h1da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_474; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1592 = 10'h1db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_475; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1593 = 10'h1dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_476; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1594 = 10'h1dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_477; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1595 = 10'h1de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_478; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1596 = 10'h1df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_479; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1597 = 10'h1e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_480; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1598 = 10'h1e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_481; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1599 = 10'h1e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_482; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1600 = 10'h1e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_483; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1601 = 10'h1e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_484; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1602 = 10'h1e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_485; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1603 = 10'h1e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_486; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1604 = 10'h1e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_487; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1605 = 10'h1e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_488; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1606 = 10'h1e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_489; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1607 = 10'h1ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_490; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1608 = 10'h1eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_491; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1609 = 10'h1ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_492; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1610 = 10'h1ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_493; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1611 = 10'h1ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_494; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1612 = 10'h1ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_495; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1613 = 10'h1f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_496; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1614 = 10'h1f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_497; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1615 = 10'h1f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_498; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1616 = 10'h1f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_499; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1617 = 10'h1f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_500; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1618 = 10'h1f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_501; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1619 = 10'h1f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_502; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1620 = 10'h1f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_503; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1621 = 10'h1f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_504; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1622 = 10'h1f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_505; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1623 = 10'h1fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_506; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1624 = 10'h1fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_507; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1625 = 10'h1fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_508; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1626 = 10'h1fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_509; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1627 = 10'h1fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_510; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1628 = 10'h1ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_511; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1629 = 10'h200 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_512; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1630 = 10'h201 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_513; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1631 = 10'h202 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_514; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1632 = 10'h203 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_515; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1633 = 10'h204 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_516; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1634 = 10'h205 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_517; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1635 = 10'h206 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_518; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1636 = 10'h207 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_519; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1637 = 10'h208 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_520; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1638 = 10'h209 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_521; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1639 = 10'h20a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_522; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1640 = 10'h20b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_523; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1641 = 10'h20c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_524; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1642 = 10'h20d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_525; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1643 = 10'h20e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_526; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1644 = 10'h20f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_527; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1645 = 10'h210 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_528; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1646 = 10'h211 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_529; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1647 = 10'h212 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_530; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1648 = 10'h213 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_531; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1649 = 10'h214 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_532; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1650 = 10'h215 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_533; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1651 = 10'h216 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_534; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1652 = 10'h217 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_535; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1653 = 10'h218 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_536; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1654 = 10'h219 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_537; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1655 = 10'h21a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_538; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1656 = 10'h21b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_539; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1657 = 10'h21c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_540; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1658 = 10'h21d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_541; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1659 = 10'h21e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_542; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1660 = 10'h21f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_543; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1661 = 10'h220 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_544; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1662 = 10'h221 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_545; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1663 = 10'h222 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_546; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1664 = 10'h223 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_547; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1665 = 10'h224 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_548; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1666 = 10'h225 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_549; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1667 = 10'h226 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_550; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1668 = 10'h227 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_551; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1669 = 10'h228 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_552; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1670 = 10'h229 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_553; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1671 = 10'h22a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_554; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1672 = 10'h22b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_555; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1673 = 10'h22c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_556; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1674 = 10'h22d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_557; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1675 = 10'h22e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_558; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1676 = 10'h22f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_559; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1677 = 10'h230 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_560; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1678 = 10'h231 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_561; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1679 = 10'h232 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_562; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1680 = 10'h233 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_563; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1681 = 10'h234 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_564; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1682 = 10'h235 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_565; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1683 = 10'h236 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_566; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1684 = 10'h237 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_567; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1685 = 10'h238 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_568; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1686 = 10'h239 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_569; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1687 = 10'h23a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_570; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1688 = 10'h23b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_571; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1689 = 10'h23c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_572; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1690 = 10'h23d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_573; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1691 = 10'h23e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_574; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1692 = 10'h23f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_575; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1693 = 10'h240 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_576; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1694 = 10'h241 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_577; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1695 = 10'h242 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_578; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1696 = 10'h243 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_579; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1697 = 10'h244 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_580; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1698 = 10'h245 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_581; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1699 = 10'h246 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_582; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1700 = 10'h247 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_583; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1701 = 10'h248 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_584; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1702 = 10'h249 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_585; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1703 = 10'h24a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_586; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1704 = 10'h24b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_587; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1705 = 10'h24c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_588; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1706 = 10'h24d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_589; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1707 = 10'h24e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_590; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1708 = 10'h24f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_591; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1709 = 10'h250 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_592; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1710 = 10'h251 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_593; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1711 = 10'h252 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_594; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1712 = 10'h253 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_595; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1713 = 10'h254 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_596; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1714 = 10'h255 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_597; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1715 = 10'h256 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_598; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1716 = 10'h257 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_599; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1717 = 10'h258 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_600; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1718 = 10'h259 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_601; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1719 = 10'h25a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_602; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1720 = 10'h25b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_603; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1721 = 10'h25c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_604; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1722 = 10'h25d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_605; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1723 = 10'h25e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_606; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1724 = 10'h25f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_607; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1725 = 10'h260 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_608; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1726 = 10'h261 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_609; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1727 = 10'h262 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_610; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1728 = 10'h263 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_611; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1729 = 10'h264 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_612; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1730 = 10'h265 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_613; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1731 = 10'h266 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_614; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1732 = 10'h267 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_615; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1733 = 10'h268 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_616; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1734 = 10'h269 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_617; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1735 = 10'h26a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_618; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1736 = 10'h26b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_619; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1737 = 10'h26c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_620; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1738 = 10'h26d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_621; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1739 = 10'h26e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_622; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1740 = 10'h26f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_623; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1741 = 10'h270 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_624; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1742 = 10'h271 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_625; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1743 = 10'h272 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_626; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1744 = 10'h273 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_627; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1745 = 10'h274 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_628; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1746 = 10'h275 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_629; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1747 = 10'h276 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_630; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1748 = 10'h277 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_631; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1749 = 10'h278 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_632; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1750 = 10'h279 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_633; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1751 = 10'h27a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_634; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1752 = 10'h27b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_635; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1753 = 10'h27c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_636; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1754 = 10'h27d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_637; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1755 = 10'h27e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_638; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1756 = 10'h27f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_639; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1757 = 10'h280 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_640; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1758 = 10'h281 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_641; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1759 = 10'h282 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_642; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1760 = 10'h283 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_643; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1761 = 10'h284 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_644; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1762 = 10'h285 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_645; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1763 = 10'h286 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_646; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1764 = 10'h287 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_647; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1765 = 10'h288 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_648; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1766 = 10'h289 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_649; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1767 = 10'h28a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_650; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1768 = 10'h28b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_651; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1769 = 10'h28c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_652; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1770 = 10'h28d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_653; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1771 = 10'h28e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_654; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1772 = 10'h28f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_655; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1773 = 10'h290 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_656; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1774 = 10'h291 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_657; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1775 = 10'h292 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_658; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1776 = 10'h293 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_659; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1777 = 10'h294 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_660; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1778 = 10'h295 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_661; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1779 = 10'h296 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_662; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1780 = 10'h297 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_663; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1781 = 10'h298 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_664; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1782 = 10'h299 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_665; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1783 = 10'h29a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_666; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1784 = 10'h29b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_667; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1785 = 10'h29c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_668; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1786 = 10'h29d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_669; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1787 = 10'h29e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_670; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1788 = 10'h29f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_671; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1789 = 10'h2a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_672; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1790 = 10'h2a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_673; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1791 = 10'h2a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_674; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1792 = 10'h2a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_675; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1793 = 10'h2a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_676; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1794 = 10'h2a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_677; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1795 = 10'h2a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_678; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1796 = 10'h2a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_679; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1797 = 10'h2a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_680; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1798 = 10'h2a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_681; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1799 = 10'h2aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_682; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1800 = 10'h2ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_683; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1801 = 10'h2ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_684; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1802 = 10'h2ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_685; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1803 = 10'h2ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_686; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1804 = 10'h2af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_687; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1805 = 10'h2b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_688; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1806 = 10'h2b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_689; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1807 = 10'h2b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_690; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1808 = 10'h2b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_691; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1809 = 10'h2b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_692; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1810 = 10'h2b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_693; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1811 = 10'h2b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_694; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1812 = 10'h2b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_695; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1813 = 10'h2b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_696; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1814 = 10'h2b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_697; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1815 = 10'h2ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_698; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1816 = 10'h2bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_699; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1817 = 10'h2bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_700; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1818 = 10'h2bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_701; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1819 = 10'h2be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_702; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1820 = 10'h2bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_703; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1821 = 10'h2c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_704; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1822 = 10'h2c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_705; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1823 = 10'h2c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_706; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1824 = 10'h2c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_707; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1825 = 10'h2c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_708; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1826 = 10'h2c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_709; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1827 = 10'h2c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_710; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1828 = 10'h2c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_711; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1829 = 10'h2c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_712; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1830 = 10'h2c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_713; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1831 = 10'h2ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_714; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1832 = 10'h2cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_715; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1833 = 10'h2cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_716; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1834 = 10'h2cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_717; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1835 = 10'h2ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_718; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1836 = 10'h2cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_719; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1837 = 10'h2d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_720; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1838 = 10'h2d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_721; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1839 = 10'h2d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_722; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1840 = 10'h2d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_723; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1841 = 10'h2d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_724; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1842 = 10'h2d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_725; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1843 = 10'h2d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_726; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1844 = 10'h2d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_727; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1845 = 10'h2d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_728; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1846 = 10'h2d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_729; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1847 = 10'h2da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_730; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1848 = 10'h2db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_731; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1849 = 10'h2dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_732; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1850 = 10'h2dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_733; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1851 = 10'h2de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_734; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1852 = 10'h2df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_735; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1853 = 10'h2e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_736; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1854 = 10'h2e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_737; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1855 = 10'h2e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_738; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1856 = 10'h2e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_739; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1857 = 10'h2e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_740; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1858 = 10'h2e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_741; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1859 = 10'h2e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_742; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1860 = 10'h2e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_743; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1861 = 10'h2e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_744; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1862 = 10'h2e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_745; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1863 = 10'h2ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_746; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1864 = 10'h2eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_747; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1865 = 10'h2ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_748; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1866 = 10'h2ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_749; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1867 = 10'h2ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_750; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1868 = 10'h2ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_751; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1869 = 10'h2f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_752; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1870 = 10'h2f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_753; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1871 = 10'h2f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_754; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1872 = 10'h2f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_755; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1873 = 10'h2f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_756; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1874 = 10'h2f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_757; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1875 = 10'h2f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_758; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1876 = 10'h2f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_759; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1877 = 10'h2f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_760; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1878 = 10'h2f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_761; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1879 = 10'h2fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_762; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1880 = 10'h2fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_763; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1881 = 10'h2fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_764; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1882 = 10'h2fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_765; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1883 = 10'h2fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_766; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1884 = 10'h2ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_767; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1885 = 10'h300 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_768; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1886 = 10'h301 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_769; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1887 = 10'h302 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_770; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1888 = 10'h303 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_771; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1889 = 10'h304 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_772; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1890 = 10'h305 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_773; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1891 = 10'h306 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_774; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1892 = 10'h307 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_775; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1893 = 10'h308 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_776; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1894 = 10'h309 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_777; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1895 = 10'h30a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_778; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1896 = 10'h30b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_779; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1897 = 10'h30c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_780; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1898 = 10'h30d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_781; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1899 = 10'h30e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_782; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1900 = 10'h30f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_783; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1901 = 10'h310 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_784; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1902 = 10'h311 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_785; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1903 = 10'h312 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_786; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1904 = 10'h313 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_787; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1905 = 10'h314 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_788; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1906 = 10'h315 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_789; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1907 = 10'h316 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_790; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1908 = 10'h317 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_791; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1909 = 10'h318 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_792; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1910 = 10'h319 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_793; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1911 = 10'h31a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_794; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1912 = 10'h31b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_795; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1913 = 10'h31c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_796; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1914 = 10'h31d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_797; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1915 = 10'h31e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_798; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1916 = 10'h31f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_799; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1917 = 10'h320 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_800; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1918 = 10'h321 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_801; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1919 = 10'h322 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_802; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1920 = 10'h323 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_803; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1921 = 10'h324 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_804; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1922 = 10'h325 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_805; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1923 = 10'h326 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_806; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1924 = 10'h327 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_807; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1925 = 10'h328 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_808; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1926 = 10'h329 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_809; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1927 = 10'h32a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_810; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1928 = 10'h32b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_811; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1929 = 10'h32c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_812; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1930 = 10'h32d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_813; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1931 = 10'h32e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_814; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1932 = 10'h32f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_815; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1933 = 10'h330 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_816; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1934 = 10'h331 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_817; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1935 = 10'h332 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_818; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1936 = 10'h333 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_819; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1937 = 10'h334 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_820; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1938 = 10'h335 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_821; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1939 = 10'h336 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_822; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1940 = 10'h337 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_823; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1941 = 10'h338 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_824; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1942 = 10'h339 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_825; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1943 = 10'h33a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_826; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1944 = 10'h33b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_827; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1945 = 10'h33c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_828; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1946 = 10'h33d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_829; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1947 = 10'h33e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_830; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1948 = 10'h33f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_831; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1949 = 10'h340 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_832; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1950 = 10'h341 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_833; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1951 = 10'h342 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_834; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1952 = 10'h343 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_835; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1953 = 10'h344 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_836; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1954 = 10'h345 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_837; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1955 = 10'h346 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_838; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1956 = 10'h347 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_839; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1957 = 10'h348 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_840; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1958 = 10'h349 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_841; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1959 = 10'h34a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_842; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1960 = 10'h34b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_843; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1961 = 10'h34c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_844; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1962 = 10'h34d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_845; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1963 = 10'h34e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_846; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1964 = 10'h34f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_847; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1965 = 10'h350 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_848; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1966 = 10'h351 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_849; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1967 = 10'h352 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_850; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1968 = 10'h353 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_851; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1969 = 10'h354 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_852; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1970 = 10'h355 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_853; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1971 = 10'h356 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_854; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1972 = 10'h357 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_855; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1973 = 10'h358 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_856; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1974 = 10'h359 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_857; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1975 = 10'h35a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_858; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1976 = 10'h35b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_859; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1977 = 10'h35c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_860; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1978 = 10'h35d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_861; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1979 = 10'h35e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_862; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1980 = 10'h35f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_863; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1981 = 10'h360 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_864; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1982 = 10'h361 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_865; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1983 = 10'h362 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_866; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1984 = 10'h363 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_867; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1985 = 10'h364 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_868; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1986 = 10'h365 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_869; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1987 = 10'h366 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_870; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1988 = 10'h367 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_871; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1989 = 10'h368 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_872; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1990 = 10'h369 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_873; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1991 = 10'h36a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_874; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1992 = 10'h36b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_875; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1993 = 10'h36c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_876; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1994 = 10'h36d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_877; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1995 = 10'h36e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_878; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1996 = 10'h36f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_879; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1997 = 10'h370 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_880; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1998 = 10'h371 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_881; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_1999 = 10'h372 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_882; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2000 = 10'h373 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_883; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2001 = 10'h374 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_884; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2002 = 10'h375 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_885; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2003 = 10'h376 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_886; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2004 = 10'h377 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_887; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2005 = 10'h378 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_888; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2006 = 10'h379 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_889; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2007 = 10'h37a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_890; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2008 = 10'h37b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_891; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2009 = 10'h37c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_892; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2010 = 10'h37d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_893; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2011 = 10'h37e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_894; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2012 = 10'h37f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_895; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2013 = 10'h380 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_896; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2014 = 10'h381 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_897; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2015 = 10'h382 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_898; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2016 = 10'h383 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_899; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2017 = 10'h384 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_900; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2018 = 10'h385 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_901; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2019 = 10'h386 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_902; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2020 = 10'h387 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_903; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2021 = 10'h388 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_904; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2022 = 10'h389 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_905; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2023 = 10'h38a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_906; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2024 = 10'h38b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_907; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2025 = 10'h38c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_908; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2026 = 10'h38d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_909; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2027 = 10'h38e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_910; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2028 = 10'h38f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_911; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2029 = 10'h390 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_912; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2030 = 10'h391 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_913; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2031 = 10'h392 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_914; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2032 = 10'h393 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_915; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2033 = 10'h394 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_916; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2034 = 10'h395 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_917; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2035 = 10'h396 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_918; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2036 = 10'h397 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_919; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2037 = 10'h398 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_920; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2038 = 10'h399 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_921; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2039 = 10'h39a == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_922; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2040 = 10'h39b == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_923; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2041 = 10'h39c == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_924; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2042 = 10'h39d == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_925; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2043 = 10'h39e == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_926; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2044 = 10'h39f == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_927; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2045 = 10'h3a0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_928; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2046 = 10'h3a1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_929; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2047 = 10'h3a2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_930; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2048 = 10'h3a3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_931; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2049 = 10'h3a4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_932; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2050 = 10'h3a5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_933; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2051 = 10'h3a6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_934; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2052 = 10'h3a7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_935; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2053 = 10'h3a8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_936; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2054 = 10'h3a9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_937; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2055 = 10'h3aa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_938; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2056 = 10'h3ab == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_939; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2057 = 10'h3ac == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_940; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2058 = 10'h3ad == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_941; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2059 = 10'h3ae == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_942; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2060 = 10'h3af == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_943; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2061 = 10'h3b0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_944; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2062 = 10'h3b1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_945; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2063 = 10'h3b2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_946; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2064 = 10'h3b3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_947; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2065 = 10'h3b4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_948; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2066 = 10'h3b5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_949; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2067 = 10'h3b6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_950; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2068 = 10'h3b7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_951; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2069 = 10'h3b8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_952; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2070 = 10'h3b9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_953; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2071 = 10'h3ba == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_954; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2072 = 10'h3bb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_955; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2073 = 10'h3bc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_956; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2074 = 10'h3bd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_957; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2075 = 10'h3be == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_958; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2076 = 10'h3bf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_959; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2077 = 10'h3c0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_960; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2078 = 10'h3c1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_961; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2079 = 10'h3c2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_962; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2080 = 10'h3c3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_963; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2081 = 10'h3c4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_964; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2082 = 10'h3c5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_965; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2083 = 10'h3c6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_966; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2084 = 10'h3c7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_967; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2085 = 10'h3c8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_968; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2086 = 10'h3c9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_969; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2087 = 10'h3ca == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_970; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2088 = 10'h3cb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_971; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2089 = 10'h3cc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_972; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2090 = 10'h3cd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_973; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2091 = 10'h3ce == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_974; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2092 = 10'h3cf == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_975; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2093 = 10'h3d0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_976; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2094 = 10'h3d1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_977; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2095 = 10'h3d2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_978; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2096 = 10'h3d3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_979; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2097 = 10'h3d4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_980; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2098 = 10'h3d5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_981; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2099 = 10'h3d6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_982; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2100 = 10'h3d7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_983; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2101 = 10'h3d8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_984; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2102 = 10'h3d9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_985; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2103 = 10'h3da == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_986; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2104 = 10'h3db == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_987; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2105 = 10'h3dc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_988; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2106 = 10'h3dd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_989; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2107 = 10'h3de == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_990; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2108 = 10'h3df == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_991; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2109 = 10'h3e0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_992; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2110 = 10'h3e1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_993; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2111 = 10'h3e2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_994; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2112 = 10'h3e3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_995; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2113 = 10'h3e4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_996; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2114 = 10'h3e5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_997; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2115 = 10'h3e6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_998; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2116 = 10'h3e7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_999; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2117 = 10'h3e8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1000; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2118 = 10'h3e9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1001; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2119 = 10'h3ea == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1002; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2120 = 10'h3eb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1003; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2121 = 10'h3ec == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1004; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2122 = 10'h3ed == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1005; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2123 = 10'h3ee == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1006; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2124 = 10'h3ef == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1007; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2125 = 10'h3f0 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1008; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2126 = 10'h3f1 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1009; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2127 = 10'h3f2 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1010; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2128 = 10'h3f3 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1011; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2129 = 10'h3f4 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1012; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2130 = 10'h3f5 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1013; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2131 = 10'h3f6 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1014; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2132 = 10'h3f7 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1015; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2133 = 10'h3f8 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1016; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2134 = 10'h3f9 == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1017; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2135 = 10'h3fa == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1018; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2136 = 10'h3fb == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1019; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2137 = 10'h3fc == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1020; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2138 = 10'h3fd == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1021; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2139 = 10'h3fe == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1022; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2140 = 10'h3ff == EXMEMALUOut[9:0] ? EXMEMB[31:0] : DMemory_1023; // @[cpu.scala 282:24 437:{37,37}]
  wire [31:0] _GEN_2141 = EXMEMop == 7'h23 ? _GEN_1117 : DMemory_0; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2142 = EXMEMop == 7'h23 ? _GEN_1118 : DMemory_1; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2143 = EXMEMop == 7'h23 ? _GEN_1119 : DMemory_2; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2144 = EXMEMop == 7'h23 ? _GEN_1120 : DMemory_3; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2145 = EXMEMop == 7'h23 ? _GEN_1121 : DMemory_4; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2146 = EXMEMop == 7'h23 ? _GEN_1122 : DMemory_5; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2147 = EXMEMop == 7'h23 ? _GEN_1123 : DMemory_6; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2148 = EXMEMop == 7'h23 ? _GEN_1124 : DMemory_7; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2149 = EXMEMop == 7'h23 ? _GEN_1125 : DMemory_8; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2150 = EXMEMop == 7'h23 ? _GEN_1126 : DMemory_9; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2151 = EXMEMop == 7'h23 ? _GEN_1127 : DMemory_10; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2152 = EXMEMop == 7'h23 ? _GEN_1128 : DMemory_11; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2153 = EXMEMop == 7'h23 ? _GEN_1129 : DMemory_12; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2154 = EXMEMop == 7'h23 ? _GEN_1130 : DMemory_13; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2155 = EXMEMop == 7'h23 ? _GEN_1131 : DMemory_14; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2156 = EXMEMop == 7'h23 ? _GEN_1132 : DMemory_15; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2157 = EXMEMop == 7'h23 ? _GEN_1133 : DMemory_16; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2158 = EXMEMop == 7'h23 ? _GEN_1134 : DMemory_17; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2159 = EXMEMop == 7'h23 ? _GEN_1135 : DMemory_18; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2160 = EXMEMop == 7'h23 ? _GEN_1136 : DMemory_19; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2161 = EXMEMop == 7'h23 ? _GEN_1137 : DMemory_20; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2162 = EXMEMop == 7'h23 ? _GEN_1138 : DMemory_21; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2163 = EXMEMop == 7'h23 ? _GEN_1139 : DMemory_22; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2164 = EXMEMop == 7'h23 ? _GEN_1140 : DMemory_23; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2165 = EXMEMop == 7'h23 ? _GEN_1141 : DMemory_24; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2166 = EXMEMop == 7'h23 ? _GEN_1142 : DMemory_25; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2167 = EXMEMop == 7'h23 ? _GEN_1143 : DMemory_26; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2168 = EXMEMop == 7'h23 ? _GEN_1144 : DMemory_27; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2169 = EXMEMop == 7'h23 ? _GEN_1145 : DMemory_28; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2170 = EXMEMop == 7'h23 ? _GEN_1146 : DMemory_29; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2171 = EXMEMop == 7'h23 ? _GEN_1147 : DMemory_30; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2172 = EXMEMop == 7'h23 ? _GEN_1148 : DMemory_31; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2173 = EXMEMop == 7'h23 ? _GEN_1149 : DMemory_32; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2174 = EXMEMop == 7'h23 ? _GEN_1150 : DMemory_33; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2175 = EXMEMop == 7'h23 ? _GEN_1151 : DMemory_34; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2176 = EXMEMop == 7'h23 ? _GEN_1152 : DMemory_35; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2177 = EXMEMop == 7'h23 ? _GEN_1153 : DMemory_36; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2178 = EXMEMop == 7'h23 ? _GEN_1154 : DMemory_37; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2179 = EXMEMop == 7'h23 ? _GEN_1155 : DMemory_38; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2180 = EXMEMop == 7'h23 ? _GEN_1156 : DMemory_39; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2181 = EXMEMop == 7'h23 ? _GEN_1157 : DMemory_40; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2182 = EXMEMop == 7'h23 ? _GEN_1158 : DMemory_41; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2183 = EXMEMop == 7'h23 ? _GEN_1159 : DMemory_42; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2184 = EXMEMop == 7'h23 ? _GEN_1160 : DMemory_43; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2185 = EXMEMop == 7'h23 ? _GEN_1161 : DMemory_44; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2186 = EXMEMop == 7'h23 ? _GEN_1162 : DMemory_45; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2187 = EXMEMop == 7'h23 ? _GEN_1163 : DMemory_46; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2188 = EXMEMop == 7'h23 ? _GEN_1164 : DMemory_47; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2189 = EXMEMop == 7'h23 ? _GEN_1165 : DMemory_48; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2190 = EXMEMop == 7'h23 ? _GEN_1166 : DMemory_49; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2191 = EXMEMop == 7'h23 ? _GEN_1167 : DMemory_50; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2192 = EXMEMop == 7'h23 ? _GEN_1168 : DMemory_51; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2193 = EXMEMop == 7'h23 ? _GEN_1169 : DMemory_52; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2194 = EXMEMop == 7'h23 ? _GEN_1170 : DMemory_53; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2195 = EXMEMop == 7'h23 ? _GEN_1171 : DMemory_54; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2196 = EXMEMop == 7'h23 ? _GEN_1172 : DMemory_55; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2197 = EXMEMop == 7'h23 ? _GEN_1173 : DMemory_56; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2198 = EXMEMop == 7'h23 ? _GEN_1174 : DMemory_57; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2199 = EXMEMop == 7'h23 ? _GEN_1175 : DMemory_58; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2200 = EXMEMop == 7'h23 ? _GEN_1176 : DMemory_59; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2201 = EXMEMop == 7'h23 ? _GEN_1177 : DMemory_60; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2202 = EXMEMop == 7'h23 ? _GEN_1178 : DMemory_61; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2203 = EXMEMop == 7'h23 ? _GEN_1179 : DMemory_62; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2204 = EXMEMop == 7'h23 ? _GEN_1180 : DMemory_63; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2205 = EXMEMop == 7'h23 ? _GEN_1181 : DMemory_64; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2206 = EXMEMop == 7'h23 ? _GEN_1182 : DMemory_65; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2207 = EXMEMop == 7'h23 ? _GEN_1183 : DMemory_66; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2208 = EXMEMop == 7'h23 ? _GEN_1184 : DMemory_67; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2209 = EXMEMop == 7'h23 ? _GEN_1185 : DMemory_68; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2210 = EXMEMop == 7'h23 ? _GEN_1186 : DMemory_69; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2211 = EXMEMop == 7'h23 ? _GEN_1187 : DMemory_70; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2212 = EXMEMop == 7'h23 ? _GEN_1188 : DMemory_71; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2213 = EXMEMop == 7'h23 ? _GEN_1189 : DMemory_72; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2214 = EXMEMop == 7'h23 ? _GEN_1190 : DMemory_73; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2215 = EXMEMop == 7'h23 ? _GEN_1191 : DMemory_74; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2216 = EXMEMop == 7'h23 ? _GEN_1192 : DMemory_75; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2217 = EXMEMop == 7'h23 ? _GEN_1193 : DMemory_76; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2218 = EXMEMop == 7'h23 ? _GEN_1194 : DMemory_77; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2219 = EXMEMop == 7'h23 ? _GEN_1195 : DMemory_78; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2220 = EXMEMop == 7'h23 ? _GEN_1196 : DMemory_79; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2221 = EXMEMop == 7'h23 ? _GEN_1197 : DMemory_80; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2222 = EXMEMop == 7'h23 ? _GEN_1198 : DMemory_81; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2223 = EXMEMop == 7'h23 ? _GEN_1199 : DMemory_82; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2224 = EXMEMop == 7'h23 ? _GEN_1200 : DMemory_83; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2225 = EXMEMop == 7'h23 ? _GEN_1201 : DMemory_84; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2226 = EXMEMop == 7'h23 ? _GEN_1202 : DMemory_85; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2227 = EXMEMop == 7'h23 ? _GEN_1203 : DMemory_86; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2228 = EXMEMop == 7'h23 ? _GEN_1204 : DMemory_87; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2229 = EXMEMop == 7'h23 ? _GEN_1205 : DMemory_88; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2230 = EXMEMop == 7'h23 ? _GEN_1206 : DMemory_89; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2231 = EXMEMop == 7'h23 ? _GEN_1207 : DMemory_90; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2232 = EXMEMop == 7'h23 ? _GEN_1208 : DMemory_91; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2233 = EXMEMop == 7'h23 ? _GEN_1209 : DMemory_92; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2234 = EXMEMop == 7'h23 ? _GEN_1210 : DMemory_93; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2235 = EXMEMop == 7'h23 ? _GEN_1211 : DMemory_94; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2236 = EXMEMop == 7'h23 ? _GEN_1212 : DMemory_95; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2237 = EXMEMop == 7'h23 ? _GEN_1213 : DMemory_96; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2238 = EXMEMop == 7'h23 ? _GEN_1214 : DMemory_97; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2239 = EXMEMop == 7'h23 ? _GEN_1215 : DMemory_98; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2240 = EXMEMop == 7'h23 ? _GEN_1216 : DMemory_99; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2241 = EXMEMop == 7'h23 ? _GEN_1217 : DMemory_100; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2242 = EXMEMop == 7'h23 ? _GEN_1218 : DMemory_101; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2243 = EXMEMop == 7'h23 ? _GEN_1219 : DMemory_102; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2244 = EXMEMop == 7'h23 ? _GEN_1220 : DMemory_103; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2245 = EXMEMop == 7'h23 ? _GEN_1221 : DMemory_104; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2246 = EXMEMop == 7'h23 ? _GEN_1222 : DMemory_105; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2247 = EXMEMop == 7'h23 ? _GEN_1223 : DMemory_106; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2248 = EXMEMop == 7'h23 ? _GEN_1224 : DMemory_107; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2249 = EXMEMop == 7'h23 ? _GEN_1225 : DMemory_108; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2250 = EXMEMop == 7'h23 ? _GEN_1226 : DMemory_109; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2251 = EXMEMop == 7'h23 ? _GEN_1227 : DMemory_110; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2252 = EXMEMop == 7'h23 ? _GEN_1228 : DMemory_111; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2253 = EXMEMop == 7'h23 ? _GEN_1229 : DMemory_112; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2254 = EXMEMop == 7'h23 ? _GEN_1230 : DMemory_113; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2255 = EXMEMop == 7'h23 ? _GEN_1231 : DMemory_114; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2256 = EXMEMop == 7'h23 ? _GEN_1232 : DMemory_115; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2257 = EXMEMop == 7'h23 ? _GEN_1233 : DMemory_116; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2258 = EXMEMop == 7'h23 ? _GEN_1234 : DMemory_117; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2259 = EXMEMop == 7'h23 ? _GEN_1235 : DMemory_118; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2260 = EXMEMop == 7'h23 ? _GEN_1236 : DMemory_119; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2261 = EXMEMop == 7'h23 ? _GEN_1237 : DMemory_120; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2262 = EXMEMop == 7'h23 ? _GEN_1238 : DMemory_121; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2263 = EXMEMop == 7'h23 ? _GEN_1239 : DMemory_122; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2264 = EXMEMop == 7'h23 ? _GEN_1240 : DMemory_123; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2265 = EXMEMop == 7'h23 ? _GEN_1241 : DMemory_124; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2266 = EXMEMop == 7'h23 ? _GEN_1242 : DMemory_125; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2267 = EXMEMop == 7'h23 ? _GEN_1243 : DMemory_126; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2268 = EXMEMop == 7'h23 ? _GEN_1244 : DMemory_127; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2269 = EXMEMop == 7'h23 ? _GEN_1245 : DMemory_128; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2270 = EXMEMop == 7'h23 ? _GEN_1246 : DMemory_129; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2271 = EXMEMop == 7'h23 ? _GEN_1247 : DMemory_130; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2272 = EXMEMop == 7'h23 ? _GEN_1248 : DMemory_131; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2273 = EXMEMop == 7'h23 ? _GEN_1249 : DMemory_132; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2274 = EXMEMop == 7'h23 ? _GEN_1250 : DMemory_133; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2275 = EXMEMop == 7'h23 ? _GEN_1251 : DMemory_134; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2276 = EXMEMop == 7'h23 ? _GEN_1252 : DMemory_135; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2277 = EXMEMop == 7'h23 ? _GEN_1253 : DMemory_136; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2278 = EXMEMop == 7'h23 ? _GEN_1254 : DMemory_137; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2279 = EXMEMop == 7'h23 ? _GEN_1255 : DMemory_138; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2280 = EXMEMop == 7'h23 ? _GEN_1256 : DMemory_139; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2281 = EXMEMop == 7'h23 ? _GEN_1257 : DMemory_140; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2282 = EXMEMop == 7'h23 ? _GEN_1258 : DMemory_141; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2283 = EXMEMop == 7'h23 ? _GEN_1259 : DMemory_142; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2284 = EXMEMop == 7'h23 ? _GEN_1260 : DMemory_143; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2285 = EXMEMop == 7'h23 ? _GEN_1261 : DMemory_144; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2286 = EXMEMop == 7'h23 ? _GEN_1262 : DMemory_145; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2287 = EXMEMop == 7'h23 ? _GEN_1263 : DMemory_146; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2288 = EXMEMop == 7'h23 ? _GEN_1264 : DMemory_147; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2289 = EXMEMop == 7'h23 ? _GEN_1265 : DMemory_148; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2290 = EXMEMop == 7'h23 ? _GEN_1266 : DMemory_149; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2291 = EXMEMop == 7'h23 ? _GEN_1267 : DMemory_150; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2292 = EXMEMop == 7'h23 ? _GEN_1268 : DMemory_151; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2293 = EXMEMop == 7'h23 ? _GEN_1269 : DMemory_152; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2294 = EXMEMop == 7'h23 ? _GEN_1270 : DMemory_153; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2295 = EXMEMop == 7'h23 ? _GEN_1271 : DMemory_154; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2296 = EXMEMop == 7'h23 ? _GEN_1272 : DMemory_155; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2297 = EXMEMop == 7'h23 ? _GEN_1273 : DMemory_156; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2298 = EXMEMop == 7'h23 ? _GEN_1274 : DMemory_157; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2299 = EXMEMop == 7'h23 ? _GEN_1275 : DMemory_158; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2300 = EXMEMop == 7'h23 ? _GEN_1276 : DMemory_159; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2301 = EXMEMop == 7'h23 ? _GEN_1277 : DMemory_160; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2302 = EXMEMop == 7'h23 ? _GEN_1278 : DMemory_161; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2303 = EXMEMop == 7'h23 ? _GEN_1279 : DMemory_162; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2304 = EXMEMop == 7'h23 ? _GEN_1280 : DMemory_163; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2305 = EXMEMop == 7'h23 ? _GEN_1281 : DMemory_164; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2306 = EXMEMop == 7'h23 ? _GEN_1282 : DMemory_165; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2307 = EXMEMop == 7'h23 ? _GEN_1283 : DMemory_166; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2308 = EXMEMop == 7'h23 ? _GEN_1284 : DMemory_167; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2309 = EXMEMop == 7'h23 ? _GEN_1285 : DMemory_168; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2310 = EXMEMop == 7'h23 ? _GEN_1286 : DMemory_169; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2311 = EXMEMop == 7'h23 ? _GEN_1287 : DMemory_170; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2312 = EXMEMop == 7'h23 ? _GEN_1288 : DMemory_171; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2313 = EXMEMop == 7'h23 ? _GEN_1289 : DMemory_172; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2314 = EXMEMop == 7'h23 ? _GEN_1290 : DMemory_173; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2315 = EXMEMop == 7'h23 ? _GEN_1291 : DMemory_174; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2316 = EXMEMop == 7'h23 ? _GEN_1292 : DMemory_175; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2317 = EXMEMop == 7'h23 ? _GEN_1293 : DMemory_176; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2318 = EXMEMop == 7'h23 ? _GEN_1294 : DMemory_177; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2319 = EXMEMop == 7'h23 ? _GEN_1295 : DMemory_178; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2320 = EXMEMop == 7'h23 ? _GEN_1296 : DMemory_179; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2321 = EXMEMop == 7'h23 ? _GEN_1297 : DMemory_180; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2322 = EXMEMop == 7'h23 ? _GEN_1298 : DMemory_181; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2323 = EXMEMop == 7'h23 ? _GEN_1299 : DMemory_182; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2324 = EXMEMop == 7'h23 ? _GEN_1300 : DMemory_183; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2325 = EXMEMop == 7'h23 ? _GEN_1301 : DMemory_184; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2326 = EXMEMop == 7'h23 ? _GEN_1302 : DMemory_185; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2327 = EXMEMop == 7'h23 ? _GEN_1303 : DMemory_186; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2328 = EXMEMop == 7'h23 ? _GEN_1304 : DMemory_187; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2329 = EXMEMop == 7'h23 ? _GEN_1305 : DMemory_188; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2330 = EXMEMop == 7'h23 ? _GEN_1306 : DMemory_189; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2331 = EXMEMop == 7'h23 ? _GEN_1307 : DMemory_190; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2332 = EXMEMop == 7'h23 ? _GEN_1308 : DMemory_191; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2333 = EXMEMop == 7'h23 ? _GEN_1309 : DMemory_192; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2334 = EXMEMop == 7'h23 ? _GEN_1310 : DMemory_193; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2335 = EXMEMop == 7'h23 ? _GEN_1311 : DMemory_194; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2336 = EXMEMop == 7'h23 ? _GEN_1312 : DMemory_195; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2337 = EXMEMop == 7'h23 ? _GEN_1313 : DMemory_196; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2338 = EXMEMop == 7'h23 ? _GEN_1314 : DMemory_197; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2339 = EXMEMop == 7'h23 ? _GEN_1315 : DMemory_198; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2340 = EXMEMop == 7'h23 ? _GEN_1316 : DMemory_199; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2341 = EXMEMop == 7'h23 ? _GEN_1317 : DMemory_200; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2342 = EXMEMop == 7'h23 ? _GEN_1318 : DMemory_201; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2343 = EXMEMop == 7'h23 ? _GEN_1319 : DMemory_202; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2344 = EXMEMop == 7'h23 ? _GEN_1320 : DMemory_203; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2345 = EXMEMop == 7'h23 ? _GEN_1321 : DMemory_204; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2346 = EXMEMop == 7'h23 ? _GEN_1322 : DMemory_205; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2347 = EXMEMop == 7'h23 ? _GEN_1323 : DMemory_206; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2348 = EXMEMop == 7'h23 ? _GEN_1324 : DMemory_207; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2349 = EXMEMop == 7'h23 ? _GEN_1325 : DMemory_208; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2350 = EXMEMop == 7'h23 ? _GEN_1326 : DMemory_209; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2351 = EXMEMop == 7'h23 ? _GEN_1327 : DMemory_210; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2352 = EXMEMop == 7'h23 ? _GEN_1328 : DMemory_211; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2353 = EXMEMop == 7'h23 ? _GEN_1329 : DMemory_212; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2354 = EXMEMop == 7'h23 ? _GEN_1330 : DMemory_213; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2355 = EXMEMop == 7'h23 ? _GEN_1331 : DMemory_214; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2356 = EXMEMop == 7'h23 ? _GEN_1332 : DMemory_215; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2357 = EXMEMop == 7'h23 ? _GEN_1333 : DMemory_216; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2358 = EXMEMop == 7'h23 ? _GEN_1334 : DMemory_217; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2359 = EXMEMop == 7'h23 ? _GEN_1335 : DMemory_218; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2360 = EXMEMop == 7'h23 ? _GEN_1336 : DMemory_219; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2361 = EXMEMop == 7'h23 ? _GEN_1337 : DMemory_220; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2362 = EXMEMop == 7'h23 ? _GEN_1338 : DMemory_221; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2363 = EXMEMop == 7'h23 ? _GEN_1339 : DMemory_222; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2364 = EXMEMop == 7'h23 ? _GEN_1340 : DMemory_223; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2365 = EXMEMop == 7'h23 ? _GEN_1341 : DMemory_224; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2366 = EXMEMop == 7'h23 ? _GEN_1342 : DMemory_225; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2367 = EXMEMop == 7'h23 ? _GEN_1343 : DMemory_226; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2368 = EXMEMop == 7'h23 ? _GEN_1344 : DMemory_227; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2369 = EXMEMop == 7'h23 ? _GEN_1345 : DMemory_228; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2370 = EXMEMop == 7'h23 ? _GEN_1346 : DMemory_229; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2371 = EXMEMop == 7'h23 ? _GEN_1347 : DMemory_230; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2372 = EXMEMop == 7'h23 ? _GEN_1348 : DMemory_231; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2373 = EXMEMop == 7'h23 ? _GEN_1349 : DMemory_232; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2374 = EXMEMop == 7'h23 ? _GEN_1350 : DMemory_233; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2375 = EXMEMop == 7'h23 ? _GEN_1351 : DMemory_234; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2376 = EXMEMop == 7'h23 ? _GEN_1352 : DMemory_235; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2377 = EXMEMop == 7'h23 ? _GEN_1353 : DMemory_236; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2378 = EXMEMop == 7'h23 ? _GEN_1354 : DMemory_237; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2379 = EXMEMop == 7'h23 ? _GEN_1355 : DMemory_238; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2380 = EXMEMop == 7'h23 ? _GEN_1356 : DMemory_239; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2381 = EXMEMop == 7'h23 ? _GEN_1357 : DMemory_240; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2382 = EXMEMop == 7'h23 ? _GEN_1358 : DMemory_241; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2383 = EXMEMop == 7'h23 ? _GEN_1359 : DMemory_242; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2384 = EXMEMop == 7'h23 ? _GEN_1360 : DMemory_243; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2385 = EXMEMop == 7'h23 ? _GEN_1361 : DMemory_244; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2386 = EXMEMop == 7'h23 ? _GEN_1362 : DMemory_245; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2387 = EXMEMop == 7'h23 ? _GEN_1363 : DMemory_246; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2388 = EXMEMop == 7'h23 ? _GEN_1364 : DMemory_247; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2389 = EXMEMop == 7'h23 ? _GEN_1365 : DMemory_248; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2390 = EXMEMop == 7'h23 ? _GEN_1366 : DMemory_249; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2391 = EXMEMop == 7'h23 ? _GEN_1367 : DMemory_250; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2392 = EXMEMop == 7'h23 ? _GEN_1368 : DMemory_251; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2393 = EXMEMop == 7'h23 ? _GEN_1369 : DMemory_252; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2394 = EXMEMop == 7'h23 ? _GEN_1370 : DMemory_253; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2395 = EXMEMop == 7'h23 ? _GEN_1371 : DMemory_254; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2396 = EXMEMop == 7'h23 ? _GEN_1372 : DMemory_255; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2397 = EXMEMop == 7'h23 ? _GEN_1373 : DMemory_256; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2398 = EXMEMop == 7'h23 ? _GEN_1374 : DMemory_257; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2399 = EXMEMop == 7'h23 ? _GEN_1375 : DMemory_258; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2400 = EXMEMop == 7'h23 ? _GEN_1376 : DMemory_259; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2401 = EXMEMop == 7'h23 ? _GEN_1377 : DMemory_260; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2402 = EXMEMop == 7'h23 ? _GEN_1378 : DMemory_261; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2403 = EXMEMop == 7'h23 ? _GEN_1379 : DMemory_262; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2404 = EXMEMop == 7'h23 ? _GEN_1380 : DMemory_263; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2405 = EXMEMop == 7'h23 ? _GEN_1381 : DMemory_264; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2406 = EXMEMop == 7'h23 ? _GEN_1382 : DMemory_265; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2407 = EXMEMop == 7'h23 ? _GEN_1383 : DMemory_266; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2408 = EXMEMop == 7'h23 ? _GEN_1384 : DMemory_267; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2409 = EXMEMop == 7'h23 ? _GEN_1385 : DMemory_268; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2410 = EXMEMop == 7'h23 ? _GEN_1386 : DMemory_269; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2411 = EXMEMop == 7'h23 ? _GEN_1387 : DMemory_270; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2412 = EXMEMop == 7'h23 ? _GEN_1388 : DMemory_271; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2413 = EXMEMop == 7'h23 ? _GEN_1389 : DMemory_272; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2414 = EXMEMop == 7'h23 ? _GEN_1390 : DMemory_273; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2415 = EXMEMop == 7'h23 ? _GEN_1391 : DMemory_274; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2416 = EXMEMop == 7'h23 ? _GEN_1392 : DMemory_275; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2417 = EXMEMop == 7'h23 ? _GEN_1393 : DMemory_276; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2418 = EXMEMop == 7'h23 ? _GEN_1394 : DMemory_277; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2419 = EXMEMop == 7'h23 ? _GEN_1395 : DMemory_278; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2420 = EXMEMop == 7'h23 ? _GEN_1396 : DMemory_279; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2421 = EXMEMop == 7'h23 ? _GEN_1397 : DMemory_280; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2422 = EXMEMop == 7'h23 ? _GEN_1398 : DMemory_281; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2423 = EXMEMop == 7'h23 ? _GEN_1399 : DMemory_282; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2424 = EXMEMop == 7'h23 ? _GEN_1400 : DMemory_283; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2425 = EXMEMop == 7'h23 ? _GEN_1401 : DMemory_284; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2426 = EXMEMop == 7'h23 ? _GEN_1402 : DMemory_285; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2427 = EXMEMop == 7'h23 ? _GEN_1403 : DMemory_286; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2428 = EXMEMop == 7'h23 ? _GEN_1404 : DMemory_287; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2429 = EXMEMop == 7'h23 ? _GEN_1405 : DMemory_288; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2430 = EXMEMop == 7'h23 ? _GEN_1406 : DMemory_289; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2431 = EXMEMop == 7'h23 ? _GEN_1407 : DMemory_290; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2432 = EXMEMop == 7'h23 ? _GEN_1408 : DMemory_291; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2433 = EXMEMop == 7'h23 ? _GEN_1409 : DMemory_292; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2434 = EXMEMop == 7'h23 ? _GEN_1410 : DMemory_293; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2435 = EXMEMop == 7'h23 ? _GEN_1411 : DMemory_294; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2436 = EXMEMop == 7'h23 ? _GEN_1412 : DMemory_295; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2437 = EXMEMop == 7'h23 ? _GEN_1413 : DMemory_296; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2438 = EXMEMop == 7'h23 ? _GEN_1414 : DMemory_297; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2439 = EXMEMop == 7'h23 ? _GEN_1415 : DMemory_298; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2440 = EXMEMop == 7'h23 ? _GEN_1416 : DMemory_299; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2441 = EXMEMop == 7'h23 ? _GEN_1417 : DMemory_300; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2442 = EXMEMop == 7'h23 ? _GEN_1418 : DMemory_301; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2443 = EXMEMop == 7'h23 ? _GEN_1419 : DMemory_302; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2444 = EXMEMop == 7'h23 ? _GEN_1420 : DMemory_303; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2445 = EXMEMop == 7'h23 ? _GEN_1421 : DMemory_304; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2446 = EXMEMop == 7'h23 ? _GEN_1422 : DMemory_305; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2447 = EXMEMop == 7'h23 ? _GEN_1423 : DMemory_306; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2448 = EXMEMop == 7'h23 ? _GEN_1424 : DMemory_307; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2449 = EXMEMop == 7'h23 ? _GEN_1425 : DMemory_308; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2450 = EXMEMop == 7'h23 ? _GEN_1426 : DMemory_309; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2451 = EXMEMop == 7'h23 ? _GEN_1427 : DMemory_310; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2452 = EXMEMop == 7'h23 ? _GEN_1428 : DMemory_311; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2453 = EXMEMop == 7'h23 ? _GEN_1429 : DMemory_312; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2454 = EXMEMop == 7'h23 ? _GEN_1430 : DMemory_313; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2455 = EXMEMop == 7'h23 ? _GEN_1431 : DMemory_314; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2456 = EXMEMop == 7'h23 ? _GEN_1432 : DMemory_315; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2457 = EXMEMop == 7'h23 ? _GEN_1433 : DMemory_316; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2458 = EXMEMop == 7'h23 ? _GEN_1434 : DMemory_317; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2459 = EXMEMop == 7'h23 ? _GEN_1435 : DMemory_318; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2460 = EXMEMop == 7'h23 ? _GEN_1436 : DMemory_319; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2461 = EXMEMop == 7'h23 ? _GEN_1437 : DMemory_320; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2462 = EXMEMop == 7'h23 ? _GEN_1438 : DMemory_321; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2463 = EXMEMop == 7'h23 ? _GEN_1439 : DMemory_322; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2464 = EXMEMop == 7'h23 ? _GEN_1440 : DMemory_323; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2465 = EXMEMop == 7'h23 ? _GEN_1441 : DMemory_324; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2466 = EXMEMop == 7'h23 ? _GEN_1442 : DMemory_325; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2467 = EXMEMop == 7'h23 ? _GEN_1443 : DMemory_326; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2468 = EXMEMop == 7'h23 ? _GEN_1444 : DMemory_327; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2469 = EXMEMop == 7'h23 ? _GEN_1445 : DMemory_328; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2470 = EXMEMop == 7'h23 ? _GEN_1446 : DMemory_329; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2471 = EXMEMop == 7'h23 ? _GEN_1447 : DMemory_330; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2472 = EXMEMop == 7'h23 ? _GEN_1448 : DMemory_331; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2473 = EXMEMop == 7'h23 ? _GEN_1449 : DMemory_332; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2474 = EXMEMop == 7'h23 ? _GEN_1450 : DMemory_333; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2475 = EXMEMop == 7'h23 ? _GEN_1451 : DMemory_334; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2476 = EXMEMop == 7'h23 ? _GEN_1452 : DMemory_335; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2477 = EXMEMop == 7'h23 ? _GEN_1453 : DMemory_336; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2478 = EXMEMop == 7'h23 ? _GEN_1454 : DMemory_337; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2479 = EXMEMop == 7'h23 ? _GEN_1455 : DMemory_338; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2480 = EXMEMop == 7'h23 ? _GEN_1456 : DMemory_339; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2481 = EXMEMop == 7'h23 ? _GEN_1457 : DMemory_340; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2482 = EXMEMop == 7'h23 ? _GEN_1458 : DMemory_341; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2483 = EXMEMop == 7'h23 ? _GEN_1459 : DMemory_342; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2484 = EXMEMop == 7'h23 ? _GEN_1460 : DMemory_343; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2485 = EXMEMop == 7'h23 ? _GEN_1461 : DMemory_344; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2486 = EXMEMop == 7'h23 ? _GEN_1462 : DMemory_345; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2487 = EXMEMop == 7'h23 ? _GEN_1463 : DMemory_346; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2488 = EXMEMop == 7'h23 ? _GEN_1464 : DMemory_347; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2489 = EXMEMop == 7'h23 ? _GEN_1465 : DMemory_348; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2490 = EXMEMop == 7'h23 ? _GEN_1466 : DMemory_349; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2491 = EXMEMop == 7'h23 ? _GEN_1467 : DMemory_350; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2492 = EXMEMop == 7'h23 ? _GEN_1468 : DMemory_351; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2493 = EXMEMop == 7'h23 ? _GEN_1469 : DMemory_352; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2494 = EXMEMop == 7'h23 ? _GEN_1470 : DMemory_353; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2495 = EXMEMop == 7'h23 ? _GEN_1471 : DMemory_354; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2496 = EXMEMop == 7'h23 ? _GEN_1472 : DMemory_355; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2497 = EXMEMop == 7'h23 ? _GEN_1473 : DMemory_356; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2498 = EXMEMop == 7'h23 ? _GEN_1474 : DMemory_357; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2499 = EXMEMop == 7'h23 ? _GEN_1475 : DMemory_358; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2500 = EXMEMop == 7'h23 ? _GEN_1476 : DMemory_359; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2501 = EXMEMop == 7'h23 ? _GEN_1477 : DMemory_360; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2502 = EXMEMop == 7'h23 ? _GEN_1478 : DMemory_361; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2503 = EXMEMop == 7'h23 ? _GEN_1479 : DMemory_362; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2504 = EXMEMop == 7'h23 ? _GEN_1480 : DMemory_363; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2505 = EXMEMop == 7'h23 ? _GEN_1481 : DMemory_364; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2506 = EXMEMop == 7'h23 ? _GEN_1482 : DMemory_365; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2507 = EXMEMop == 7'h23 ? _GEN_1483 : DMemory_366; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2508 = EXMEMop == 7'h23 ? _GEN_1484 : DMemory_367; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2509 = EXMEMop == 7'h23 ? _GEN_1485 : DMemory_368; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2510 = EXMEMop == 7'h23 ? _GEN_1486 : DMemory_369; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2511 = EXMEMop == 7'h23 ? _GEN_1487 : DMemory_370; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2512 = EXMEMop == 7'h23 ? _GEN_1488 : DMemory_371; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2513 = EXMEMop == 7'h23 ? _GEN_1489 : DMemory_372; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2514 = EXMEMop == 7'h23 ? _GEN_1490 : DMemory_373; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2515 = EXMEMop == 7'h23 ? _GEN_1491 : DMemory_374; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2516 = EXMEMop == 7'h23 ? _GEN_1492 : DMemory_375; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2517 = EXMEMop == 7'h23 ? _GEN_1493 : DMemory_376; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2518 = EXMEMop == 7'h23 ? _GEN_1494 : DMemory_377; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2519 = EXMEMop == 7'h23 ? _GEN_1495 : DMemory_378; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2520 = EXMEMop == 7'h23 ? _GEN_1496 : DMemory_379; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2521 = EXMEMop == 7'h23 ? _GEN_1497 : DMemory_380; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2522 = EXMEMop == 7'h23 ? _GEN_1498 : DMemory_381; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2523 = EXMEMop == 7'h23 ? _GEN_1499 : DMemory_382; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2524 = EXMEMop == 7'h23 ? _GEN_1500 : DMemory_383; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2525 = EXMEMop == 7'h23 ? _GEN_1501 : DMemory_384; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2526 = EXMEMop == 7'h23 ? _GEN_1502 : DMemory_385; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2527 = EXMEMop == 7'h23 ? _GEN_1503 : DMemory_386; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2528 = EXMEMop == 7'h23 ? _GEN_1504 : DMemory_387; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2529 = EXMEMop == 7'h23 ? _GEN_1505 : DMemory_388; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2530 = EXMEMop == 7'h23 ? _GEN_1506 : DMemory_389; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2531 = EXMEMop == 7'h23 ? _GEN_1507 : DMemory_390; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2532 = EXMEMop == 7'h23 ? _GEN_1508 : DMemory_391; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2533 = EXMEMop == 7'h23 ? _GEN_1509 : DMemory_392; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2534 = EXMEMop == 7'h23 ? _GEN_1510 : DMemory_393; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2535 = EXMEMop == 7'h23 ? _GEN_1511 : DMemory_394; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2536 = EXMEMop == 7'h23 ? _GEN_1512 : DMemory_395; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2537 = EXMEMop == 7'h23 ? _GEN_1513 : DMemory_396; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2538 = EXMEMop == 7'h23 ? _GEN_1514 : DMemory_397; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2539 = EXMEMop == 7'h23 ? _GEN_1515 : DMemory_398; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2540 = EXMEMop == 7'h23 ? _GEN_1516 : DMemory_399; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2541 = EXMEMop == 7'h23 ? _GEN_1517 : DMemory_400; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2542 = EXMEMop == 7'h23 ? _GEN_1518 : DMemory_401; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2543 = EXMEMop == 7'h23 ? _GEN_1519 : DMemory_402; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2544 = EXMEMop == 7'h23 ? _GEN_1520 : DMemory_403; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2545 = EXMEMop == 7'h23 ? _GEN_1521 : DMemory_404; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2546 = EXMEMop == 7'h23 ? _GEN_1522 : DMemory_405; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2547 = EXMEMop == 7'h23 ? _GEN_1523 : DMemory_406; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2548 = EXMEMop == 7'h23 ? _GEN_1524 : DMemory_407; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2549 = EXMEMop == 7'h23 ? _GEN_1525 : DMemory_408; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2550 = EXMEMop == 7'h23 ? _GEN_1526 : DMemory_409; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2551 = EXMEMop == 7'h23 ? _GEN_1527 : DMemory_410; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2552 = EXMEMop == 7'h23 ? _GEN_1528 : DMemory_411; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2553 = EXMEMop == 7'h23 ? _GEN_1529 : DMemory_412; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2554 = EXMEMop == 7'h23 ? _GEN_1530 : DMemory_413; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2555 = EXMEMop == 7'h23 ? _GEN_1531 : DMemory_414; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2556 = EXMEMop == 7'h23 ? _GEN_1532 : DMemory_415; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2557 = EXMEMop == 7'h23 ? _GEN_1533 : DMemory_416; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2558 = EXMEMop == 7'h23 ? _GEN_1534 : DMemory_417; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2559 = EXMEMop == 7'h23 ? _GEN_1535 : DMemory_418; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2560 = EXMEMop == 7'h23 ? _GEN_1536 : DMemory_419; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2561 = EXMEMop == 7'h23 ? _GEN_1537 : DMemory_420; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2562 = EXMEMop == 7'h23 ? _GEN_1538 : DMemory_421; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2563 = EXMEMop == 7'h23 ? _GEN_1539 : DMemory_422; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2564 = EXMEMop == 7'h23 ? _GEN_1540 : DMemory_423; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2565 = EXMEMop == 7'h23 ? _GEN_1541 : DMemory_424; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2566 = EXMEMop == 7'h23 ? _GEN_1542 : DMemory_425; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2567 = EXMEMop == 7'h23 ? _GEN_1543 : DMemory_426; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2568 = EXMEMop == 7'h23 ? _GEN_1544 : DMemory_427; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2569 = EXMEMop == 7'h23 ? _GEN_1545 : DMemory_428; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2570 = EXMEMop == 7'h23 ? _GEN_1546 : DMemory_429; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2571 = EXMEMop == 7'h23 ? _GEN_1547 : DMemory_430; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2572 = EXMEMop == 7'h23 ? _GEN_1548 : DMemory_431; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2573 = EXMEMop == 7'h23 ? _GEN_1549 : DMemory_432; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2574 = EXMEMop == 7'h23 ? _GEN_1550 : DMemory_433; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2575 = EXMEMop == 7'h23 ? _GEN_1551 : DMemory_434; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2576 = EXMEMop == 7'h23 ? _GEN_1552 : DMemory_435; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2577 = EXMEMop == 7'h23 ? _GEN_1553 : DMemory_436; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2578 = EXMEMop == 7'h23 ? _GEN_1554 : DMemory_437; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2579 = EXMEMop == 7'h23 ? _GEN_1555 : DMemory_438; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2580 = EXMEMop == 7'h23 ? _GEN_1556 : DMemory_439; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2581 = EXMEMop == 7'h23 ? _GEN_1557 : DMemory_440; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2582 = EXMEMop == 7'h23 ? _GEN_1558 : DMemory_441; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2583 = EXMEMop == 7'h23 ? _GEN_1559 : DMemory_442; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2584 = EXMEMop == 7'h23 ? _GEN_1560 : DMemory_443; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2585 = EXMEMop == 7'h23 ? _GEN_1561 : DMemory_444; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2586 = EXMEMop == 7'h23 ? _GEN_1562 : DMemory_445; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2587 = EXMEMop == 7'h23 ? _GEN_1563 : DMemory_446; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2588 = EXMEMop == 7'h23 ? _GEN_1564 : DMemory_447; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2589 = EXMEMop == 7'h23 ? _GEN_1565 : DMemory_448; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2590 = EXMEMop == 7'h23 ? _GEN_1566 : DMemory_449; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2591 = EXMEMop == 7'h23 ? _GEN_1567 : DMemory_450; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2592 = EXMEMop == 7'h23 ? _GEN_1568 : DMemory_451; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2593 = EXMEMop == 7'h23 ? _GEN_1569 : DMemory_452; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2594 = EXMEMop == 7'h23 ? _GEN_1570 : DMemory_453; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2595 = EXMEMop == 7'h23 ? _GEN_1571 : DMemory_454; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2596 = EXMEMop == 7'h23 ? _GEN_1572 : DMemory_455; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2597 = EXMEMop == 7'h23 ? _GEN_1573 : DMemory_456; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2598 = EXMEMop == 7'h23 ? _GEN_1574 : DMemory_457; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2599 = EXMEMop == 7'h23 ? _GEN_1575 : DMemory_458; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2600 = EXMEMop == 7'h23 ? _GEN_1576 : DMemory_459; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2601 = EXMEMop == 7'h23 ? _GEN_1577 : DMemory_460; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2602 = EXMEMop == 7'h23 ? _GEN_1578 : DMemory_461; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2603 = EXMEMop == 7'h23 ? _GEN_1579 : DMemory_462; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2604 = EXMEMop == 7'h23 ? _GEN_1580 : DMemory_463; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2605 = EXMEMop == 7'h23 ? _GEN_1581 : DMemory_464; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2606 = EXMEMop == 7'h23 ? _GEN_1582 : DMemory_465; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2607 = EXMEMop == 7'h23 ? _GEN_1583 : DMemory_466; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2608 = EXMEMop == 7'h23 ? _GEN_1584 : DMemory_467; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2609 = EXMEMop == 7'h23 ? _GEN_1585 : DMemory_468; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2610 = EXMEMop == 7'h23 ? _GEN_1586 : DMemory_469; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2611 = EXMEMop == 7'h23 ? _GEN_1587 : DMemory_470; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2612 = EXMEMop == 7'h23 ? _GEN_1588 : DMemory_471; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2613 = EXMEMop == 7'h23 ? _GEN_1589 : DMemory_472; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2614 = EXMEMop == 7'h23 ? _GEN_1590 : DMemory_473; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2615 = EXMEMop == 7'h23 ? _GEN_1591 : DMemory_474; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2616 = EXMEMop == 7'h23 ? _GEN_1592 : DMemory_475; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2617 = EXMEMop == 7'h23 ? _GEN_1593 : DMemory_476; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2618 = EXMEMop == 7'h23 ? _GEN_1594 : DMemory_477; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2619 = EXMEMop == 7'h23 ? _GEN_1595 : DMemory_478; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2620 = EXMEMop == 7'h23 ? _GEN_1596 : DMemory_479; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2621 = EXMEMop == 7'h23 ? _GEN_1597 : DMemory_480; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2622 = EXMEMop == 7'h23 ? _GEN_1598 : DMemory_481; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2623 = EXMEMop == 7'h23 ? _GEN_1599 : DMemory_482; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2624 = EXMEMop == 7'h23 ? _GEN_1600 : DMemory_483; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2625 = EXMEMop == 7'h23 ? _GEN_1601 : DMemory_484; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2626 = EXMEMop == 7'h23 ? _GEN_1602 : DMemory_485; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2627 = EXMEMop == 7'h23 ? _GEN_1603 : DMemory_486; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2628 = EXMEMop == 7'h23 ? _GEN_1604 : DMemory_487; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2629 = EXMEMop == 7'h23 ? _GEN_1605 : DMemory_488; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2630 = EXMEMop == 7'h23 ? _GEN_1606 : DMemory_489; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2631 = EXMEMop == 7'h23 ? _GEN_1607 : DMemory_490; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2632 = EXMEMop == 7'h23 ? _GEN_1608 : DMemory_491; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2633 = EXMEMop == 7'h23 ? _GEN_1609 : DMemory_492; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2634 = EXMEMop == 7'h23 ? _GEN_1610 : DMemory_493; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2635 = EXMEMop == 7'h23 ? _GEN_1611 : DMemory_494; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2636 = EXMEMop == 7'h23 ? _GEN_1612 : DMemory_495; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2637 = EXMEMop == 7'h23 ? _GEN_1613 : DMemory_496; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2638 = EXMEMop == 7'h23 ? _GEN_1614 : DMemory_497; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2639 = EXMEMop == 7'h23 ? _GEN_1615 : DMemory_498; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2640 = EXMEMop == 7'h23 ? _GEN_1616 : DMemory_499; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2641 = EXMEMop == 7'h23 ? _GEN_1617 : DMemory_500; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2642 = EXMEMop == 7'h23 ? _GEN_1618 : DMemory_501; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2643 = EXMEMop == 7'h23 ? _GEN_1619 : DMemory_502; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2644 = EXMEMop == 7'h23 ? _GEN_1620 : DMemory_503; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2645 = EXMEMop == 7'h23 ? _GEN_1621 : DMemory_504; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2646 = EXMEMop == 7'h23 ? _GEN_1622 : DMemory_505; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2647 = EXMEMop == 7'h23 ? _GEN_1623 : DMemory_506; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2648 = EXMEMop == 7'h23 ? _GEN_1624 : DMemory_507; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2649 = EXMEMop == 7'h23 ? _GEN_1625 : DMemory_508; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2650 = EXMEMop == 7'h23 ? _GEN_1626 : DMemory_509; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2651 = EXMEMop == 7'h23 ? _GEN_1627 : DMemory_510; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2652 = EXMEMop == 7'h23 ? _GEN_1628 : DMemory_511; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2653 = EXMEMop == 7'h23 ? _GEN_1629 : DMemory_512; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2654 = EXMEMop == 7'h23 ? _GEN_1630 : DMemory_513; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2655 = EXMEMop == 7'h23 ? _GEN_1631 : DMemory_514; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2656 = EXMEMop == 7'h23 ? _GEN_1632 : DMemory_515; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2657 = EXMEMop == 7'h23 ? _GEN_1633 : DMemory_516; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2658 = EXMEMop == 7'h23 ? _GEN_1634 : DMemory_517; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2659 = EXMEMop == 7'h23 ? _GEN_1635 : DMemory_518; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2660 = EXMEMop == 7'h23 ? _GEN_1636 : DMemory_519; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2661 = EXMEMop == 7'h23 ? _GEN_1637 : DMemory_520; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2662 = EXMEMop == 7'h23 ? _GEN_1638 : DMemory_521; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2663 = EXMEMop == 7'h23 ? _GEN_1639 : DMemory_522; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2664 = EXMEMop == 7'h23 ? _GEN_1640 : DMemory_523; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2665 = EXMEMop == 7'h23 ? _GEN_1641 : DMemory_524; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2666 = EXMEMop == 7'h23 ? _GEN_1642 : DMemory_525; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2667 = EXMEMop == 7'h23 ? _GEN_1643 : DMemory_526; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2668 = EXMEMop == 7'h23 ? _GEN_1644 : DMemory_527; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2669 = EXMEMop == 7'h23 ? _GEN_1645 : DMemory_528; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2670 = EXMEMop == 7'h23 ? _GEN_1646 : DMemory_529; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2671 = EXMEMop == 7'h23 ? _GEN_1647 : DMemory_530; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2672 = EXMEMop == 7'h23 ? _GEN_1648 : DMemory_531; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2673 = EXMEMop == 7'h23 ? _GEN_1649 : DMemory_532; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2674 = EXMEMop == 7'h23 ? _GEN_1650 : DMemory_533; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2675 = EXMEMop == 7'h23 ? _GEN_1651 : DMemory_534; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2676 = EXMEMop == 7'h23 ? _GEN_1652 : DMemory_535; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2677 = EXMEMop == 7'h23 ? _GEN_1653 : DMemory_536; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2678 = EXMEMop == 7'h23 ? _GEN_1654 : DMemory_537; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2679 = EXMEMop == 7'h23 ? _GEN_1655 : DMemory_538; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2680 = EXMEMop == 7'h23 ? _GEN_1656 : DMemory_539; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2681 = EXMEMop == 7'h23 ? _GEN_1657 : DMemory_540; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2682 = EXMEMop == 7'h23 ? _GEN_1658 : DMemory_541; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2683 = EXMEMop == 7'h23 ? _GEN_1659 : DMemory_542; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2684 = EXMEMop == 7'h23 ? _GEN_1660 : DMemory_543; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2685 = EXMEMop == 7'h23 ? _GEN_1661 : DMemory_544; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2686 = EXMEMop == 7'h23 ? _GEN_1662 : DMemory_545; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2687 = EXMEMop == 7'h23 ? _GEN_1663 : DMemory_546; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2688 = EXMEMop == 7'h23 ? _GEN_1664 : DMemory_547; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2689 = EXMEMop == 7'h23 ? _GEN_1665 : DMemory_548; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2690 = EXMEMop == 7'h23 ? _GEN_1666 : DMemory_549; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2691 = EXMEMop == 7'h23 ? _GEN_1667 : DMemory_550; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2692 = EXMEMop == 7'h23 ? _GEN_1668 : DMemory_551; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2693 = EXMEMop == 7'h23 ? _GEN_1669 : DMemory_552; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2694 = EXMEMop == 7'h23 ? _GEN_1670 : DMemory_553; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2695 = EXMEMop == 7'h23 ? _GEN_1671 : DMemory_554; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2696 = EXMEMop == 7'h23 ? _GEN_1672 : DMemory_555; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2697 = EXMEMop == 7'h23 ? _GEN_1673 : DMemory_556; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2698 = EXMEMop == 7'h23 ? _GEN_1674 : DMemory_557; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2699 = EXMEMop == 7'h23 ? _GEN_1675 : DMemory_558; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2700 = EXMEMop == 7'h23 ? _GEN_1676 : DMemory_559; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2701 = EXMEMop == 7'h23 ? _GEN_1677 : DMemory_560; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2702 = EXMEMop == 7'h23 ? _GEN_1678 : DMemory_561; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2703 = EXMEMop == 7'h23 ? _GEN_1679 : DMemory_562; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2704 = EXMEMop == 7'h23 ? _GEN_1680 : DMemory_563; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2705 = EXMEMop == 7'h23 ? _GEN_1681 : DMemory_564; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2706 = EXMEMop == 7'h23 ? _GEN_1682 : DMemory_565; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2707 = EXMEMop == 7'h23 ? _GEN_1683 : DMemory_566; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2708 = EXMEMop == 7'h23 ? _GEN_1684 : DMemory_567; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2709 = EXMEMop == 7'h23 ? _GEN_1685 : DMemory_568; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2710 = EXMEMop == 7'h23 ? _GEN_1686 : DMemory_569; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2711 = EXMEMop == 7'h23 ? _GEN_1687 : DMemory_570; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2712 = EXMEMop == 7'h23 ? _GEN_1688 : DMemory_571; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2713 = EXMEMop == 7'h23 ? _GEN_1689 : DMemory_572; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2714 = EXMEMop == 7'h23 ? _GEN_1690 : DMemory_573; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2715 = EXMEMop == 7'h23 ? _GEN_1691 : DMemory_574; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2716 = EXMEMop == 7'h23 ? _GEN_1692 : DMemory_575; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2717 = EXMEMop == 7'h23 ? _GEN_1693 : DMemory_576; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2718 = EXMEMop == 7'h23 ? _GEN_1694 : DMemory_577; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2719 = EXMEMop == 7'h23 ? _GEN_1695 : DMemory_578; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2720 = EXMEMop == 7'h23 ? _GEN_1696 : DMemory_579; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2721 = EXMEMop == 7'h23 ? _GEN_1697 : DMemory_580; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2722 = EXMEMop == 7'h23 ? _GEN_1698 : DMemory_581; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2723 = EXMEMop == 7'h23 ? _GEN_1699 : DMemory_582; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2724 = EXMEMop == 7'h23 ? _GEN_1700 : DMemory_583; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2725 = EXMEMop == 7'h23 ? _GEN_1701 : DMemory_584; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2726 = EXMEMop == 7'h23 ? _GEN_1702 : DMemory_585; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2727 = EXMEMop == 7'h23 ? _GEN_1703 : DMemory_586; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2728 = EXMEMop == 7'h23 ? _GEN_1704 : DMemory_587; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2729 = EXMEMop == 7'h23 ? _GEN_1705 : DMemory_588; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2730 = EXMEMop == 7'h23 ? _GEN_1706 : DMemory_589; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2731 = EXMEMop == 7'h23 ? _GEN_1707 : DMemory_590; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2732 = EXMEMop == 7'h23 ? _GEN_1708 : DMemory_591; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2733 = EXMEMop == 7'h23 ? _GEN_1709 : DMemory_592; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2734 = EXMEMop == 7'h23 ? _GEN_1710 : DMemory_593; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2735 = EXMEMop == 7'h23 ? _GEN_1711 : DMemory_594; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2736 = EXMEMop == 7'h23 ? _GEN_1712 : DMemory_595; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2737 = EXMEMop == 7'h23 ? _GEN_1713 : DMemory_596; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2738 = EXMEMop == 7'h23 ? _GEN_1714 : DMemory_597; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2739 = EXMEMop == 7'h23 ? _GEN_1715 : DMemory_598; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2740 = EXMEMop == 7'h23 ? _GEN_1716 : DMemory_599; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2741 = EXMEMop == 7'h23 ? _GEN_1717 : DMemory_600; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2742 = EXMEMop == 7'h23 ? _GEN_1718 : DMemory_601; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2743 = EXMEMop == 7'h23 ? _GEN_1719 : DMemory_602; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2744 = EXMEMop == 7'h23 ? _GEN_1720 : DMemory_603; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2745 = EXMEMop == 7'h23 ? _GEN_1721 : DMemory_604; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2746 = EXMEMop == 7'h23 ? _GEN_1722 : DMemory_605; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2747 = EXMEMop == 7'h23 ? _GEN_1723 : DMemory_606; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2748 = EXMEMop == 7'h23 ? _GEN_1724 : DMemory_607; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2749 = EXMEMop == 7'h23 ? _GEN_1725 : DMemory_608; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2750 = EXMEMop == 7'h23 ? _GEN_1726 : DMemory_609; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2751 = EXMEMop == 7'h23 ? _GEN_1727 : DMemory_610; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2752 = EXMEMop == 7'h23 ? _GEN_1728 : DMemory_611; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2753 = EXMEMop == 7'h23 ? _GEN_1729 : DMemory_612; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2754 = EXMEMop == 7'h23 ? _GEN_1730 : DMemory_613; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2755 = EXMEMop == 7'h23 ? _GEN_1731 : DMemory_614; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2756 = EXMEMop == 7'h23 ? _GEN_1732 : DMemory_615; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2757 = EXMEMop == 7'h23 ? _GEN_1733 : DMemory_616; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2758 = EXMEMop == 7'h23 ? _GEN_1734 : DMemory_617; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2759 = EXMEMop == 7'h23 ? _GEN_1735 : DMemory_618; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2760 = EXMEMop == 7'h23 ? _GEN_1736 : DMemory_619; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2761 = EXMEMop == 7'h23 ? _GEN_1737 : DMemory_620; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2762 = EXMEMop == 7'h23 ? _GEN_1738 : DMemory_621; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2763 = EXMEMop == 7'h23 ? _GEN_1739 : DMemory_622; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2764 = EXMEMop == 7'h23 ? _GEN_1740 : DMemory_623; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2765 = EXMEMop == 7'h23 ? _GEN_1741 : DMemory_624; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2766 = EXMEMop == 7'h23 ? _GEN_1742 : DMemory_625; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2767 = EXMEMop == 7'h23 ? _GEN_1743 : DMemory_626; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2768 = EXMEMop == 7'h23 ? _GEN_1744 : DMemory_627; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2769 = EXMEMop == 7'h23 ? _GEN_1745 : DMemory_628; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2770 = EXMEMop == 7'h23 ? _GEN_1746 : DMemory_629; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2771 = EXMEMop == 7'h23 ? _GEN_1747 : DMemory_630; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2772 = EXMEMop == 7'h23 ? _GEN_1748 : DMemory_631; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2773 = EXMEMop == 7'h23 ? _GEN_1749 : DMemory_632; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2774 = EXMEMop == 7'h23 ? _GEN_1750 : DMemory_633; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2775 = EXMEMop == 7'h23 ? _GEN_1751 : DMemory_634; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2776 = EXMEMop == 7'h23 ? _GEN_1752 : DMemory_635; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2777 = EXMEMop == 7'h23 ? _GEN_1753 : DMemory_636; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2778 = EXMEMop == 7'h23 ? _GEN_1754 : DMemory_637; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2779 = EXMEMop == 7'h23 ? _GEN_1755 : DMemory_638; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2780 = EXMEMop == 7'h23 ? _GEN_1756 : DMemory_639; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2781 = EXMEMop == 7'h23 ? _GEN_1757 : DMemory_640; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2782 = EXMEMop == 7'h23 ? _GEN_1758 : DMemory_641; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2783 = EXMEMop == 7'h23 ? _GEN_1759 : DMemory_642; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2784 = EXMEMop == 7'h23 ? _GEN_1760 : DMemory_643; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2785 = EXMEMop == 7'h23 ? _GEN_1761 : DMemory_644; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2786 = EXMEMop == 7'h23 ? _GEN_1762 : DMemory_645; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2787 = EXMEMop == 7'h23 ? _GEN_1763 : DMemory_646; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2788 = EXMEMop == 7'h23 ? _GEN_1764 : DMemory_647; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2789 = EXMEMop == 7'h23 ? _GEN_1765 : DMemory_648; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2790 = EXMEMop == 7'h23 ? _GEN_1766 : DMemory_649; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2791 = EXMEMop == 7'h23 ? _GEN_1767 : DMemory_650; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2792 = EXMEMop == 7'h23 ? _GEN_1768 : DMemory_651; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2793 = EXMEMop == 7'h23 ? _GEN_1769 : DMemory_652; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2794 = EXMEMop == 7'h23 ? _GEN_1770 : DMemory_653; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2795 = EXMEMop == 7'h23 ? _GEN_1771 : DMemory_654; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2796 = EXMEMop == 7'h23 ? _GEN_1772 : DMemory_655; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2797 = EXMEMop == 7'h23 ? _GEN_1773 : DMemory_656; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2798 = EXMEMop == 7'h23 ? _GEN_1774 : DMemory_657; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2799 = EXMEMop == 7'h23 ? _GEN_1775 : DMemory_658; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2800 = EXMEMop == 7'h23 ? _GEN_1776 : DMemory_659; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2801 = EXMEMop == 7'h23 ? _GEN_1777 : DMemory_660; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2802 = EXMEMop == 7'h23 ? _GEN_1778 : DMemory_661; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2803 = EXMEMop == 7'h23 ? _GEN_1779 : DMemory_662; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2804 = EXMEMop == 7'h23 ? _GEN_1780 : DMemory_663; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2805 = EXMEMop == 7'h23 ? _GEN_1781 : DMemory_664; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2806 = EXMEMop == 7'h23 ? _GEN_1782 : DMemory_665; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2807 = EXMEMop == 7'h23 ? _GEN_1783 : DMemory_666; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2808 = EXMEMop == 7'h23 ? _GEN_1784 : DMemory_667; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2809 = EXMEMop == 7'h23 ? _GEN_1785 : DMemory_668; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2810 = EXMEMop == 7'h23 ? _GEN_1786 : DMemory_669; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2811 = EXMEMop == 7'h23 ? _GEN_1787 : DMemory_670; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2812 = EXMEMop == 7'h23 ? _GEN_1788 : DMemory_671; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2813 = EXMEMop == 7'h23 ? _GEN_1789 : DMemory_672; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2814 = EXMEMop == 7'h23 ? _GEN_1790 : DMemory_673; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2815 = EXMEMop == 7'h23 ? _GEN_1791 : DMemory_674; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2816 = EXMEMop == 7'h23 ? _GEN_1792 : DMemory_675; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2817 = EXMEMop == 7'h23 ? _GEN_1793 : DMemory_676; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2818 = EXMEMop == 7'h23 ? _GEN_1794 : DMemory_677; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2819 = EXMEMop == 7'h23 ? _GEN_1795 : DMemory_678; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2820 = EXMEMop == 7'h23 ? _GEN_1796 : DMemory_679; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2821 = EXMEMop == 7'h23 ? _GEN_1797 : DMemory_680; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2822 = EXMEMop == 7'h23 ? _GEN_1798 : DMemory_681; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2823 = EXMEMop == 7'h23 ? _GEN_1799 : DMemory_682; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2824 = EXMEMop == 7'h23 ? _GEN_1800 : DMemory_683; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2825 = EXMEMop == 7'h23 ? _GEN_1801 : DMemory_684; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2826 = EXMEMop == 7'h23 ? _GEN_1802 : DMemory_685; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2827 = EXMEMop == 7'h23 ? _GEN_1803 : DMemory_686; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2828 = EXMEMop == 7'h23 ? _GEN_1804 : DMemory_687; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2829 = EXMEMop == 7'h23 ? _GEN_1805 : DMemory_688; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2830 = EXMEMop == 7'h23 ? _GEN_1806 : DMemory_689; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2831 = EXMEMop == 7'h23 ? _GEN_1807 : DMemory_690; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2832 = EXMEMop == 7'h23 ? _GEN_1808 : DMemory_691; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2833 = EXMEMop == 7'h23 ? _GEN_1809 : DMemory_692; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2834 = EXMEMop == 7'h23 ? _GEN_1810 : DMemory_693; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2835 = EXMEMop == 7'h23 ? _GEN_1811 : DMemory_694; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2836 = EXMEMop == 7'h23 ? _GEN_1812 : DMemory_695; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2837 = EXMEMop == 7'h23 ? _GEN_1813 : DMemory_696; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2838 = EXMEMop == 7'h23 ? _GEN_1814 : DMemory_697; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2839 = EXMEMop == 7'h23 ? _GEN_1815 : DMemory_698; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2840 = EXMEMop == 7'h23 ? _GEN_1816 : DMemory_699; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2841 = EXMEMop == 7'h23 ? _GEN_1817 : DMemory_700; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2842 = EXMEMop == 7'h23 ? _GEN_1818 : DMemory_701; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2843 = EXMEMop == 7'h23 ? _GEN_1819 : DMemory_702; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2844 = EXMEMop == 7'h23 ? _GEN_1820 : DMemory_703; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2845 = EXMEMop == 7'h23 ? _GEN_1821 : DMemory_704; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2846 = EXMEMop == 7'h23 ? _GEN_1822 : DMemory_705; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2847 = EXMEMop == 7'h23 ? _GEN_1823 : DMemory_706; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2848 = EXMEMop == 7'h23 ? _GEN_1824 : DMemory_707; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2849 = EXMEMop == 7'h23 ? _GEN_1825 : DMemory_708; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2850 = EXMEMop == 7'h23 ? _GEN_1826 : DMemory_709; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2851 = EXMEMop == 7'h23 ? _GEN_1827 : DMemory_710; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2852 = EXMEMop == 7'h23 ? _GEN_1828 : DMemory_711; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2853 = EXMEMop == 7'h23 ? _GEN_1829 : DMemory_712; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2854 = EXMEMop == 7'h23 ? _GEN_1830 : DMemory_713; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2855 = EXMEMop == 7'h23 ? _GEN_1831 : DMemory_714; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2856 = EXMEMop == 7'h23 ? _GEN_1832 : DMemory_715; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2857 = EXMEMop == 7'h23 ? _GEN_1833 : DMemory_716; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2858 = EXMEMop == 7'h23 ? _GEN_1834 : DMemory_717; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2859 = EXMEMop == 7'h23 ? _GEN_1835 : DMemory_718; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2860 = EXMEMop == 7'h23 ? _GEN_1836 : DMemory_719; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2861 = EXMEMop == 7'h23 ? _GEN_1837 : DMemory_720; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2862 = EXMEMop == 7'h23 ? _GEN_1838 : DMemory_721; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2863 = EXMEMop == 7'h23 ? _GEN_1839 : DMemory_722; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2864 = EXMEMop == 7'h23 ? _GEN_1840 : DMemory_723; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2865 = EXMEMop == 7'h23 ? _GEN_1841 : DMemory_724; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2866 = EXMEMop == 7'h23 ? _GEN_1842 : DMemory_725; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2867 = EXMEMop == 7'h23 ? _GEN_1843 : DMemory_726; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2868 = EXMEMop == 7'h23 ? _GEN_1844 : DMemory_727; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2869 = EXMEMop == 7'h23 ? _GEN_1845 : DMemory_728; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2870 = EXMEMop == 7'h23 ? _GEN_1846 : DMemory_729; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2871 = EXMEMop == 7'h23 ? _GEN_1847 : DMemory_730; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2872 = EXMEMop == 7'h23 ? _GEN_1848 : DMemory_731; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2873 = EXMEMop == 7'h23 ? _GEN_1849 : DMemory_732; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2874 = EXMEMop == 7'h23 ? _GEN_1850 : DMemory_733; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2875 = EXMEMop == 7'h23 ? _GEN_1851 : DMemory_734; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2876 = EXMEMop == 7'h23 ? _GEN_1852 : DMemory_735; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2877 = EXMEMop == 7'h23 ? _GEN_1853 : DMemory_736; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2878 = EXMEMop == 7'h23 ? _GEN_1854 : DMemory_737; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2879 = EXMEMop == 7'h23 ? _GEN_1855 : DMemory_738; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2880 = EXMEMop == 7'h23 ? _GEN_1856 : DMemory_739; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2881 = EXMEMop == 7'h23 ? _GEN_1857 : DMemory_740; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2882 = EXMEMop == 7'h23 ? _GEN_1858 : DMemory_741; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2883 = EXMEMop == 7'h23 ? _GEN_1859 : DMemory_742; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2884 = EXMEMop == 7'h23 ? _GEN_1860 : DMemory_743; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2885 = EXMEMop == 7'h23 ? _GEN_1861 : DMemory_744; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2886 = EXMEMop == 7'h23 ? _GEN_1862 : DMemory_745; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2887 = EXMEMop == 7'h23 ? _GEN_1863 : DMemory_746; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2888 = EXMEMop == 7'h23 ? _GEN_1864 : DMemory_747; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2889 = EXMEMop == 7'h23 ? _GEN_1865 : DMemory_748; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2890 = EXMEMop == 7'h23 ? _GEN_1866 : DMemory_749; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2891 = EXMEMop == 7'h23 ? _GEN_1867 : DMemory_750; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2892 = EXMEMop == 7'h23 ? _GEN_1868 : DMemory_751; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2893 = EXMEMop == 7'h23 ? _GEN_1869 : DMemory_752; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2894 = EXMEMop == 7'h23 ? _GEN_1870 : DMemory_753; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2895 = EXMEMop == 7'h23 ? _GEN_1871 : DMemory_754; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2896 = EXMEMop == 7'h23 ? _GEN_1872 : DMemory_755; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2897 = EXMEMop == 7'h23 ? _GEN_1873 : DMemory_756; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2898 = EXMEMop == 7'h23 ? _GEN_1874 : DMemory_757; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2899 = EXMEMop == 7'h23 ? _GEN_1875 : DMemory_758; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2900 = EXMEMop == 7'h23 ? _GEN_1876 : DMemory_759; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2901 = EXMEMop == 7'h23 ? _GEN_1877 : DMemory_760; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2902 = EXMEMop == 7'h23 ? _GEN_1878 : DMemory_761; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2903 = EXMEMop == 7'h23 ? _GEN_1879 : DMemory_762; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2904 = EXMEMop == 7'h23 ? _GEN_1880 : DMemory_763; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2905 = EXMEMop == 7'h23 ? _GEN_1881 : DMemory_764; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2906 = EXMEMop == 7'h23 ? _GEN_1882 : DMemory_765; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2907 = EXMEMop == 7'h23 ? _GEN_1883 : DMemory_766; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2908 = EXMEMop == 7'h23 ? _GEN_1884 : DMemory_767; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2909 = EXMEMop == 7'h23 ? _GEN_1885 : DMemory_768; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2910 = EXMEMop == 7'h23 ? _GEN_1886 : DMemory_769; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2911 = EXMEMop == 7'h23 ? _GEN_1887 : DMemory_770; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2912 = EXMEMop == 7'h23 ? _GEN_1888 : DMemory_771; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2913 = EXMEMop == 7'h23 ? _GEN_1889 : DMemory_772; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2914 = EXMEMop == 7'h23 ? _GEN_1890 : DMemory_773; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2915 = EXMEMop == 7'h23 ? _GEN_1891 : DMemory_774; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2916 = EXMEMop == 7'h23 ? _GEN_1892 : DMemory_775; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2917 = EXMEMop == 7'h23 ? _GEN_1893 : DMemory_776; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2918 = EXMEMop == 7'h23 ? _GEN_1894 : DMemory_777; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2919 = EXMEMop == 7'h23 ? _GEN_1895 : DMemory_778; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2920 = EXMEMop == 7'h23 ? _GEN_1896 : DMemory_779; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2921 = EXMEMop == 7'h23 ? _GEN_1897 : DMemory_780; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2922 = EXMEMop == 7'h23 ? _GEN_1898 : DMemory_781; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2923 = EXMEMop == 7'h23 ? _GEN_1899 : DMemory_782; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2924 = EXMEMop == 7'h23 ? _GEN_1900 : DMemory_783; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2925 = EXMEMop == 7'h23 ? _GEN_1901 : DMemory_784; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2926 = EXMEMop == 7'h23 ? _GEN_1902 : DMemory_785; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2927 = EXMEMop == 7'h23 ? _GEN_1903 : DMemory_786; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2928 = EXMEMop == 7'h23 ? _GEN_1904 : DMemory_787; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2929 = EXMEMop == 7'h23 ? _GEN_1905 : DMemory_788; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2930 = EXMEMop == 7'h23 ? _GEN_1906 : DMemory_789; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2931 = EXMEMop == 7'h23 ? _GEN_1907 : DMemory_790; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2932 = EXMEMop == 7'h23 ? _GEN_1908 : DMemory_791; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2933 = EXMEMop == 7'h23 ? _GEN_1909 : DMemory_792; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2934 = EXMEMop == 7'h23 ? _GEN_1910 : DMemory_793; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2935 = EXMEMop == 7'h23 ? _GEN_1911 : DMemory_794; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2936 = EXMEMop == 7'h23 ? _GEN_1912 : DMemory_795; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2937 = EXMEMop == 7'h23 ? _GEN_1913 : DMemory_796; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2938 = EXMEMop == 7'h23 ? _GEN_1914 : DMemory_797; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2939 = EXMEMop == 7'h23 ? _GEN_1915 : DMemory_798; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2940 = EXMEMop == 7'h23 ? _GEN_1916 : DMemory_799; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2941 = EXMEMop == 7'h23 ? _GEN_1917 : DMemory_800; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2942 = EXMEMop == 7'h23 ? _GEN_1918 : DMemory_801; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2943 = EXMEMop == 7'h23 ? _GEN_1919 : DMemory_802; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2944 = EXMEMop == 7'h23 ? _GEN_1920 : DMemory_803; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2945 = EXMEMop == 7'h23 ? _GEN_1921 : DMemory_804; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2946 = EXMEMop == 7'h23 ? _GEN_1922 : DMemory_805; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2947 = EXMEMop == 7'h23 ? _GEN_1923 : DMemory_806; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2948 = EXMEMop == 7'h23 ? _GEN_1924 : DMemory_807; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2949 = EXMEMop == 7'h23 ? _GEN_1925 : DMemory_808; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2950 = EXMEMop == 7'h23 ? _GEN_1926 : DMemory_809; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2951 = EXMEMop == 7'h23 ? _GEN_1927 : DMemory_810; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2952 = EXMEMop == 7'h23 ? _GEN_1928 : DMemory_811; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2953 = EXMEMop == 7'h23 ? _GEN_1929 : DMemory_812; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2954 = EXMEMop == 7'h23 ? _GEN_1930 : DMemory_813; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2955 = EXMEMop == 7'h23 ? _GEN_1931 : DMemory_814; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2956 = EXMEMop == 7'h23 ? _GEN_1932 : DMemory_815; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2957 = EXMEMop == 7'h23 ? _GEN_1933 : DMemory_816; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2958 = EXMEMop == 7'h23 ? _GEN_1934 : DMemory_817; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2959 = EXMEMop == 7'h23 ? _GEN_1935 : DMemory_818; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2960 = EXMEMop == 7'h23 ? _GEN_1936 : DMemory_819; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2961 = EXMEMop == 7'h23 ? _GEN_1937 : DMemory_820; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2962 = EXMEMop == 7'h23 ? _GEN_1938 : DMemory_821; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2963 = EXMEMop == 7'h23 ? _GEN_1939 : DMemory_822; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2964 = EXMEMop == 7'h23 ? _GEN_1940 : DMemory_823; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2965 = EXMEMop == 7'h23 ? _GEN_1941 : DMemory_824; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2966 = EXMEMop == 7'h23 ? _GEN_1942 : DMemory_825; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2967 = EXMEMop == 7'h23 ? _GEN_1943 : DMemory_826; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2968 = EXMEMop == 7'h23 ? _GEN_1944 : DMemory_827; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2969 = EXMEMop == 7'h23 ? _GEN_1945 : DMemory_828; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2970 = EXMEMop == 7'h23 ? _GEN_1946 : DMemory_829; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2971 = EXMEMop == 7'h23 ? _GEN_1947 : DMemory_830; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2972 = EXMEMop == 7'h23 ? _GEN_1948 : DMemory_831; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2973 = EXMEMop == 7'h23 ? _GEN_1949 : DMemory_832; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2974 = EXMEMop == 7'h23 ? _GEN_1950 : DMemory_833; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2975 = EXMEMop == 7'h23 ? _GEN_1951 : DMemory_834; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2976 = EXMEMop == 7'h23 ? _GEN_1952 : DMemory_835; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2977 = EXMEMop == 7'h23 ? _GEN_1953 : DMemory_836; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2978 = EXMEMop == 7'h23 ? _GEN_1954 : DMemory_837; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2979 = EXMEMop == 7'h23 ? _GEN_1955 : DMemory_838; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2980 = EXMEMop == 7'h23 ? _GEN_1956 : DMemory_839; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2981 = EXMEMop == 7'h23 ? _GEN_1957 : DMemory_840; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2982 = EXMEMop == 7'h23 ? _GEN_1958 : DMemory_841; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2983 = EXMEMop == 7'h23 ? _GEN_1959 : DMemory_842; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2984 = EXMEMop == 7'h23 ? _GEN_1960 : DMemory_843; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2985 = EXMEMop == 7'h23 ? _GEN_1961 : DMemory_844; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2986 = EXMEMop == 7'h23 ? _GEN_1962 : DMemory_845; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2987 = EXMEMop == 7'h23 ? _GEN_1963 : DMemory_846; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2988 = EXMEMop == 7'h23 ? _GEN_1964 : DMemory_847; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2989 = EXMEMop == 7'h23 ? _GEN_1965 : DMemory_848; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2990 = EXMEMop == 7'h23 ? _GEN_1966 : DMemory_849; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2991 = EXMEMop == 7'h23 ? _GEN_1967 : DMemory_850; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2992 = EXMEMop == 7'h23 ? _GEN_1968 : DMemory_851; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2993 = EXMEMop == 7'h23 ? _GEN_1969 : DMemory_852; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2994 = EXMEMop == 7'h23 ? _GEN_1970 : DMemory_853; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2995 = EXMEMop == 7'h23 ? _GEN_1971 : DMemory_854; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2996 = EXMEMop == 7'h23 ? _GEN_1972 : DMemory_855; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2997 = EXMEMop == 7'h23 ? _GEN_1973 : DMemory_856; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2998 = EXMEMop == 7'h23 ? _GEN_1974 : DMemory_857; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_2999 = EXMEMop == 7'h23 ? _GEN_1975 : DMemory_858; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3000 = EXMEMop == 7'h23 ? _GEN_1976 : DMemory_859; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3001 = EXMEMop == 7'h23 ? _GEN_1977 : DMemory_860; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3002 = EXMEMop == 7'h23 ? _GEN_1978 : DMemory_861; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3003 = EXMEMop == 7'h23 ? _GEN_1979 : DMemory_862; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3004 = EXMEMop == 7'h23 ? _GEN_1980 : DMemory_863; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3005 = EXMEMop == 7'h23 ? _GEN_1981 : DMemory_864; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3006 = EXMEMop == 7'h23 ? _GEN_1982 : DMemory_865; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3007 = EXMEMop == 7'h23 ? _GEN_1983 : DMemory_866; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3008 = EXMEMop == 7'h23 ? _GEN_1984 : DMemory_867; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3009 = EXMEMop == 7'h23 ? _GEN_1985 : DMemory_868; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3010 = EXMEMop == 7'h23 ? _GEN_1986 : DMemory_869; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3011 = EXMEMop == 7'h23 ? _GEN_1987 : DMemory_870; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3012 = EXMEMop == 7'h23 ? _GEN_1988 : DMemory_871; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3013 = EXMEMop == 7'h23 ? _GEN_1989 : DMemory_872; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3014 = EXMEMop == 7'h23 ? _GEN_1990 : DMemory_873; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3015 = EXMEMop == 7'h23 ? _GEN_1991 : DMemory_874; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3016 = EXMEMop == 7'h23 ? _GEN_1992 : DMemory_875; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3017 = EXMEMop == 7'h23 ? _GEN_1993 : DMemory_876; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3018 = EXMEMop == 7'h23 ? _GEN_1994 : DMemory_877; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3019 = EXMEMop == 7'h23 ? _GEN_1995 : DMemory_878; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3020 = EXMEMop == 7'h23 ? _GEN_1996 : DMemory_879; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3021 = EXMEMop == 7'h23 ? _GEN_1997 : DMemory_880; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3022 = EXMEMop == 7'h23 ? _GEN_1998 : DMemory_881; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3023 = EXMEMop == 7'h23 ? _GEN_1999 : DMemory_882; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3024 = EXMEMop == 7'h23 ? _GEN_2000 : DMemory_883; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3025 = EXMEMop == 7'h23 ? _GEN_2001 : DMemory_884; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3026 = EXMEMop == 7'h23 ? _GEN_2002 : DMemory_885; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3027 = EXMEMop == 7'h23 ? _GEN_2003 : DMemory_886; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3028 = EXMEMop == 7'h23 ? _GEN_2004 : DMemory_887; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3029 = EXMEMop == 7'h23 ? _GEN_2005 : DMemory_888; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3030 = EXMEMop == 7'h23 ? _GEN_2006 : DMemory_889; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3031 = EXMEMop == 7'h23 ? _GEN_2007 : DMemory_890; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3032 = EXMEMop == 7'h23 ? _GEN_2008 : DMemory_891; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3033 = EXMEMop == 7'h23 ? _GEN_2009 : DMemory_892; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3034 = EXMEMop == 7'h23 ? _GEN_2010 : DMemory_893; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3035 = EXMEMop == 7'h23 ? _GEN_2011 : DMemory_894; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3036 = EXMEMop == 7'h23 ? _GEN_2012 : DMemory_895; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3037 = EXMEMop == 7'h23 ? _GEN_2013 : DMemory_896; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3038 = EXMEMop == 7'h23 ? _GEN_2014 : DMemory_897; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3039 = EXMEMop == 7'h23 ? _GEN_2015 : DMemory_898; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3040 = EXMEMop == 7'h23 ? _GEN_2016 : DMemory_899; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3041 = EXMEMop == 7'h23 ? _GEN_2017 : DMemory_900; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3042 = EXMEMop == 7'h23 ? _GEN_2018 : DMemory_901; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3043 = EXMEMop == 7'h23 ? _GEN_2019 : DMemory_902; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3044 = EXMEMop == 7'h23 ? _GEN_2020 : DMemory_903; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3045 = EXMEMop == 7'h23 ? _GEN_2021 : DMemory_904; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3046 = EXMEMop == 7'h23 ? _GEN_2022 : DMemory_905; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3047 = EXMEMop == 7'h23 ? _GEN_2023 : DMemory_906; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3048 = EXMEMop == 7'h23 ? _GEN_2024 : DMemory_907; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3049 = EXMEMop == 7'h23 ? _GEN_2025 : DMemory_908; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3050 = EXMEMop == 7'h23 ? _GEN_2026 : DMemory_909; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3051 = EXMEMop == 7'h23 ? _GEN_2027 : DMemory_910; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3052 = EXMEMop == 7'h23 ? _GEN_2028 : DMemory_911; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3053 = EXMEMop == 7'h23 ? _GEN_2029 : DMemory_912; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3054 = EXMEMop == 7'h23 ? _GEN_2030 : DMemory_913; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3055 = EXMEMop == 7'h23 ? _GEN_2031 : DMemory_914; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3056 = EXMEMop == 7'h23 ? _GEN_2032 : DMemory_915; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3057 = EXMEMop == 7'h23 ? _GEN_2033 : DMemory_916; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3058 = EXMEMop == 7'h23 ? _GEN_2034 : DMemory_917; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3059 = EXMEMop == 7'h23 ? _GEN_2035 : DMemory_918; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3060 = EXMEMop == 7'h23 ? _GEN_2036 : DMemory_919; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3061 = EXMEMop == 7'h23 ? _GEN_2037 : DMemory_920; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3062 = EXMEMop == 7'h23 ? _GEN_2038 : DMemory_921; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3063 = EXMEMop == 7'h23 ? _GEN_2039 : DMemory_922; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3064 = EXMEMop == 7'h23 ? _GEN_2040 : DMemory_923; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3065 = EXMEMop == 7'h23 ? _GEN_2041 : DMemory_924; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3066 = EXMEMop == 7'h23 ? _GEN_2042 : DMemory_925; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3067 = EXMEMop == 7'h23 ? _GEN_2043 : DMemory_926; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3068 = EXMEMop == 7'h23 ? _GEN_2044 : DMemory_927; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3069 = EXMEMop == 7'h23 ? _GEN_2045 : DMemory_928; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3070 = EXMEMop == 7'h23 ? _GEN_2046 : DMemory_929; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3071 = EXMEMop == 7'h23 ? _GEN_2047 : DMemory_930; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3072 = EXMEMop == 7'h23 ? _GEN_2048 : DMemory_931; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3073 = EXMEMop == 7'h23 ? _GEN_2049 : DMemory_932; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3074 = EXMEMop == 7'h23 ? _GEN_2050 : DMemory_933; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3075 = EXMEMop == 7'h23 ? _GEN_2051 : DMemory_934; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3076 = EXMEMop == 7'h23 ? _GEN_2052 : DMemory_935; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3077 = EXMEMop == 7'h23 ? _GEN_2053 : DMemory_936; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3078 = EXMEMop == 7'h23 ? _GEN_2054 : DMemory_937; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3079 = EXMEMop == 7'h23 ? _GEN_2055 : DMemory_938; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3080 = EXMEMop == 7'h23 ? _GEN_2056 : DMemory_939; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3081 = EXMEMop == 7'h23 ? _GEN_2057 : DMemory_940; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3082 = EXMEMop == 7'h23 ? _GEN_2058 : DMemory_941; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3083 = EXMEMop == 7'h23 ? _GEN_2059 : DMemory_942; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3084 = EXMEMop == 7'h23 ? _GEN_2060 : DMemory_943; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3085 = EXMEMop == 7'h23 ? _GEN_2061 : DMemory_944; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3086 = EXMEMop == 7'h23 ? _GEN_2062 : DMemory_945; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3087 = EXMEMop == 7'h23 ? _GEN_2063 : DMemory_946; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3088 = EXMEMop == 7'h23 ? _GEN_2064 : DMemory_947; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3089 = EXMEMop == 7'h23 ? _GEN_2065 : DMemory_948; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3090 = EXMEMop == 7'h23 ? _GEN_2066 : DMemory_949; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3091 = EXMEMop == 7'h23 ? _GEN_2067 : DMemory_950; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3092 = EXMEMop == 7'h23 ? _GEN_2068 : DMemory_951; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3093 = EXMEMop == 7'h23 ? _GEN_2069 : DMemory_952; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3094 = EXMEMop == 7'h23 ? _GEN_2070 : DMemory_953; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3095 = EXMEMop == 7'h23 ? _GEN_2071 : DMemory_954; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3096 = EXMEMop == 7'h23 ? _GEN_2072 : DMemory_955; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3097 = EXMEMop == 7'h23 ? _GEN_2073 : DMemory_956; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3098 = EXMEMop == 7'h23 ? _GEN_2074 : DMemory_957; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3099 = EXMEMop == 7'h23 ? _GEN_2075 : DMemory_958; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3100 = EXMEMop == 7'h23 ? _GEN_2076 : DMemory_959; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3101 = EXMEMop == 7'h23 ? _GEN_2077 : DMemory_960; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3102 = EXMEMop == 7'h23 ? _GEN_2078 : DMemory_961; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3103 = EXMEMop == 7'h23 ? _GEN_2079 : DMemory_962; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3104 = EXMEMop == 7'h23 ? _GEN_2080 : DMemory_963; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3105 = EXMEMop == 7'h23 ? _GEN_2081 : DMemory_964; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3106 = EXMEMop == 7'h23 ? _GEN_2082 : DMemory_965; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3107 = EXMEMop == 7'h23 ? _GEN_2083 : DMemory_966; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3108 = EXMEMop == 7'h23 ? _GEN_2084 : DMemory_967; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3109 = EXMEMop == 7'h23 ? _GEN_2085 : DMemory_968; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3110 = EXMEMop == 7'h23 ? _GEN_2086 : DMemory_969; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3111 = EXMEMop == 7'h23 ? _GEN_2087 : DMemory_970; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3112 = EXMEMop == 7'h23 ? _GEN_2088 : DMemory_971; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3113 = EXMEMop == 7'h23 ? _GEN_2089 : DMemory_972; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3114 = EXMEMop == 7'h23 ? _GEN_2090 : DMemory_973; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3115 = EXMEMop == 7'h23 ? _GEN_2091 : DMemory_974; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3116 = EXMEMop == 7'h23 ? _GEN_2092 : DMemory_975; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3117 = EXMEMop == 7'h23 ? _GEN_2093 : DMemory_976; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3118 = EXMEMop == 7'h23 ? _GEN_2094 : DMemory_977; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3119 = EXMEMop == 7'h23 ? _GEN_2095 : DMemory_978; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3120 = EXMEMop == 7'h23 ? _GEN_2096 : DMemory_979; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3121 = EXMEMop == 7'h23 ? _GEN_2097 : DMemory_980; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3122 = EXMEMop == 7'h23 ? _GEN_2098 : DMemory_981; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3123 = EXMEMop == 7'h23 ? _GEN_2099 : DMemory_982; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3124 = EXMEMop == 7'h23 ? _GEN_2100 : DMemory_983; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3125 = EXMEMop == 7'h23 ? _GEN_2101 : DMemory_984; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3126 = EXMEMop == 7'h23 ? _GEN_2102 : DMemory_985; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3127 = EXMEMop == 7'h23 ? _GEN_2103 : DMemory_986; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3128 = EXMEMop == 7'h23 ? _GEN_2104 : DMemory_987; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3129 = EXMEMop == 7'h23 ? _GEN_2105 : DMemory_988; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3130 = EXMEMop == 7'h23 ? _GEN_2106 : DMemory_989; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3131 = EXMEMop == 7'h23 ? _GEN_2107 : DMemory_990; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3132 = EXMEMop == 7'h23 ? _GEN_2108 : DMemory_991; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3133 = EXMEMop == 7'h23 ? _GEN_2109 : DMemory_992; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3134 = EXMEMop == 7'h23 ? _GEN_2110 : DMemory_993; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3135 = EXMEMop == 7'h23 ? _GEN_2111 : DMemory_994; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3136 = EXMEMop == 7'h23 ? _GEN_2112 : DMemory_995; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3137 = EXMEMop == 7'h23 ? _GEN_2113 : DMemory_996; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3138 = EXMEMop == 7'h23 ? _GEN_2114 : DMemory_997; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3139 = EXMEMop == 7'h23 ? _GEN_2115 : DMemory_998; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3140 = EXMEMop == 7'h23 ? _GEN_2116 : DMemory_999; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3141 = EXMEMop == 7'h23 ? _GEN_2117 : DMemory_1000; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3142 = EXMEMop == 7'h23 ? _GEN_2118 : DMemory_1001; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3143 = EXMEMop == 7'h23 ? _GEN_2119 : DMemory_1002; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3144 = EXMEMop == 7'h23 ? _GEN_2120 : DMemory_1003; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3145 = EXMEMop == 7'h23 ? _GEN_2121 : DMemory_1004; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3146 = EXMEMop == 7'h23 ? _GEN_2122 : DMemory_1005; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3147 = EXMEMop == 7'h23 ? _GEN_2123 : DMemory_1006; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3148 = EXMEMop == 7'h23 ? _GEN_2124 : DMemory_1007; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3149 = EXMEMop == 7'h23 ? _GEN_2125 : DMemory_1008; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3150 = EXMEMop == 7'h23 ? _GEN_2126 : DMemory_1009; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3151 = EXMEMop == 7'h23 ? _GEN_2127 : DMemory_1010; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3152 = EXMEMop == 7'h23 ? _GEN_2128 : DMemory_1011; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3153 = EXMEMop == 7'h23 ? _GEN_2129 : DMemory_1012; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3154 = EXMEMop == 7'h23 ? _GEN_2130 : DMemory_1013; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3155 = EXMEMop == 7'h23 ? _GEN_2131 : DMemory_1014; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3156 = EXMEMop == 7'h23 ? _GEN_2132 : DMemory_1015; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3157 = EXMEMop == 7'h23 ? _GEN_2133 : DMemory_1016; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3158 = EXMEMop == 7'h23 ? _GEN_2134 : DMemory_1017; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3159 = EXMEMop == 7'h23 ? _GEN_2135 : DMemory_1018; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3160 = EXMEMop == 7'h23 ? _GEN_2136 : DMemory_1019; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3161 = EXMEMop == 7'h23 ? _GEN_2137 : DMemory_1020; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3162 = EXMEMop == 7'h23 ? _GEN_2138 : DMemory_1021; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3163 = EXMEMop == 7'h23 ? _GEN_2139 : DMemory_1022; // @[cpu.scala 282:24 436:32]
  wire [31:0] _GEN_3164 = EXMEMop == 7'h23 ? _GEN_2140 : DMemory_1023; // @[cpu.scala 282:24 436:32]
  ControlUnit ControlUnit ( // @[cpu.scala 293:20]
    .clock(ControlUnit_clock),
    .reset(ControlUnit_reset),
    .io_reset(ControlUnit_io_reset),
    .io_insns_0(ControlUnit_io_insns_0),
    .io_insns_1(ControlUnit_io_insns_1),
    .io_PC(ControlUnit_io_PC),
    .io_nPC(ControlUnit_io_nPC),
    .io_insn(ControlUnit_io_insn)
  );
  assign io_rvfi_regs_0 = Regs_0; // @[cpu.scala 453:16]
  assign io_rvfi_regs_1 = Regs_1; // @[cpu.scala 453:16]
  assign io_rvfi_regs_2 = Regs_2; // @[cpu.scala 453:16]
  assign io_rvfi_regs_3 = Regs_3; // @[cpu.scala 453:16]
  assign io_rvfi_regs_4 = Regs_4; // @[cpu.scala 453:16]
  assign io_rvfi_regs_5 = Regs_5; // @[cpu.scala 453:16]
  assign io_rvfi_regs_6 = Regs_6; // @[cpu.scala 453:16]
  assign io_rvfi_regs_7 = Regs_7; // @[cpu.scala 453:16]
  assign io_rvfi_regs_8 = Regs_8; // @[cpu.scala 453:16]
  assign io_rvfi_regs_9 = Regs_9; // @[cpu.scala 453:16]
  assign io_rvfi_regs_10 = Regs_10; // @[cpu.scala 453:16]
  assign io_rvfi_regs_11 = Regs_11; // @[cpu.scala 453:16]
  assign io_rvfi_regs_12 = Regs_12; // @[cpu.scala 453:16]
  assign io_rvfi_regs_13 = Regs_13; // @[cpu.scala 453:16]
  assign io_rvfi_regs_14 = Regs_14; // @[cpu.scala 453:16]
  assign io_rvfi_regs_15 = Regs_15; // @[cpu.scala 453:16]
  assign io_rvfi_regs_16 = Regs_16; // @[cpu.scala 453:16]
  assign io_rvfi_regs_17 = Regs_17; // @[cpu.scala 453:16]
  assign io_rvfi_regs_18 = Regs_18; // @[cpu.scala 453:16]
  assign io_rvfi_regs_19 = Regs_19; // @[cpu.scala 453:16]
  assign io_rvfi_regs_20 = Regs_20; // @[cpu.scala 453:16]
  assign io_rvfi_regs_21 = Regs_21; // @[cpu.scala 453:16]
  assign io_rvfi_regs_22 = Regs_22; // @[cpu.scala 453:16]
  assign io_rvfi_regs_23 = Regs_23; // @[cpu.scala 453:16]
  assign io_rvfi_regs_24 = Regs_24; // @[cpu.scala 453:16]
  assign io_rvfi_regs_25 = Regs_25; // @[cpu.scala 453:16]
  assign io_rvfi_regs_26 = Regs_26; // @[cpu.scala 453:16]
  assign io_rvfi_regs_27 = Regs_27; // @[cpu.scala 453:16]
  assign io_rvfi_regs_28 = Regs_28; // @[cpu.scala 453:16]
  assign io_rvfi_regs_29 = Regs_29; // @[cpu.scala 453:16]
  assign io_rvfi_regs_30 = Regs_30; // @[cpu.scala 453:16]
  assign io_rvfi_regs_31 = Regs_31; // @[cpu.scala 453:16]
  assign ControlUnit_clock = clock;
  assign ControlUnit_reset = reset;
  assign ControlUnit_io_reset = io_rvfi_rst; // @[cpu.scala 296:14]
  assign ControlUnit_io_insns_0 = IMemory_0; // @[cpu.scala 295:14]
  assign ControlUnit_io_insns_1 = IMemory_1; // @[cpu.scala 295:14]
  assign ControlUnit_io_PC = PC; // @[cpu.scala 294:11]
  always @(posedge clock) begin
    if (reset) begin // @[cpu.scala 277:19]
      PC <= 64'h0; // @[cpu.scala 277:19]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (~stall) begin // @[cpu.scala 353:27]
        if (~takeBranch) begin // @[cpu.scala 354:34]
          PC <= ControlUnit_io_nPC; // @[cpu.scala 358:12]
        end else begin
          PC <= branchTarget; // @[cpu.scala 374:12]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_0 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h0 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_0 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_1 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h1 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_1 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_2 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h2 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_2 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_3 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h3 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_3 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_4 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h4 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_4 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_5 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h5 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_5 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_6 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h6 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_6 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_7 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h7 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_7 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_8 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h8 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_8 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_9 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h9 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_9 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_10 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'ha == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_10 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_11 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'hb == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_11 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_12 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'hc == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_12 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_13 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'hd == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_13 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_14 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'he == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_14 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_15 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'hf == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_15 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_16 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h10 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_16 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_17 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h11 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_17 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_18 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h12 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_18 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_19 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h13 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_19 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_20 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h14 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_20 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_21 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h15 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_21 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_22 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h16 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_22 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_23 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h17 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_23 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_24 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h18 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_24 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_25 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h19 == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_25 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_26 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h1a == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_26 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_27 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h1b == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_27 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_28 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h1c == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_28 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_29 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h1d == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_29 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_30 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h1e == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_30 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (reset) begin // @[cpu.scala 278:21]
      Regs_31 <= 64'h0; // @[cpu.scala 278:21]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if ((_bypassAFromWB_T_4 | _bypassAFromWB_T_3) & MEMWBrd != 5'h0) begin // @[cpu.scala 446:74]
        if (5'h1f == MEMWBrd) begin // @[cpu.scala 447:21]
          Regs_31 <= MEMWBValue; // @[cpu.scala 447:21]
        end
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (~stall) begin // @[cpu.scala 353:27]
        if (bypassAFromEX) begin // @[cpu.scala 380:27]
          IDEXA <= _A_T_1; // @[cpu.scala 382:11]
        end else if (bypassAFromMEM) begin // @[cpu.scala 383:34]
          IDEXA <= EXMEMALUOut; // @[cpu.scala 385:11]
        end else begin
          IDEXA <= _GEN_37;
        end
      end else begin
        IDEXA <= 64'h0;
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (~stall) begin // @[cpu.scala 353:27]
        if (bypassBFromEX) begin // @[cpu.scala 393:27]
          IDEXB <= _B_T_1; // @[cpu.scala 395:11]
        end else if (bypassBFromMEM) begin // @[cpu.scala 396:34]
          IDEXB <= EXMEMALUOut; // @[cpu.scala 398:11]
        end else begin
          IDEXB <= _GEN_75;
        end
      end else begin
        IDEXB <= 64'h0;
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      EXMEMB <= IDEXB; // @[cpu.scala 429:12]
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (_stall_T_9) begin // @[cpu.scala 414:25]
        EXMEMALUOut <= _EXMEMALUOut_T_6; // @[cpu.scala 415:19]
      end else if (IDEXop == 7'h23) begin // @[cpu.scala 416:31]
        EXMEMALUOut <= _EXMEMALUOut_T_15; // @[cpu.scala 417:19]
      end else if (_bypassAFromEX_T_3) begin // @[cpu.scala 421:34]
        EXMEMALUOut <= _A_T_1; // @[cpu.scala 424:19]
      end
    end
    if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (_bypassAFromMEM_T_3) begin // @[cpu.scala 432:29]
        MEMWBValue <= EXMEMALUOut; // @[cpu.scala 433:18]
      end else if (_stall_T) begin // @[cpu.scala 434:32]
        MEMWBValue <= {{32'd0}, _GEN_1116}; // @[cpu.scala 435:18]
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_0 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_0 <= _GEN_2141;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1 <= _GEN_2142;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_2 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_2 <= _GEN_2143;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_3 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_3 <= _GEN_2144;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_4 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_4 <= _GEN_2145;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_5 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_5 <= _GEN_2146;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_6 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_6 <= _GEN_2147;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_7 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_7 <= _GEN_2148;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_8 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_8 <= _GEN_2149;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_9 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_9 <= _GEN_2150;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_10 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_10 <= _GEN_2151;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_11 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_11 <= _GEN_2152;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_12 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_12 <= _GEN_2153;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_13 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_13 <= _GEN_2154;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_14 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_14 <= _GEN_2155;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_15 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_15 <= _GEN_2156;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_16 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_16 <= _GEN_2157;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_17 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_17 <= _GEN_2158;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_18 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_18 <= _GEN_2159;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_19 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_19 <= _GEN_2160;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_20 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_20 <= _GEN_2161;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_21 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_21 <= _GEN_2162;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_22 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_22 <= _GEN_2163;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_23 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_23 <= _GEN_2164;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_24 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_24 <= _GEN_2165;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_25 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_25 <= _GEN_2166;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_26 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_26 <= _GEN_2167;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_27 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_27 <= _GEN_2168;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_28 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_28 <= _GEN_2169;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_29 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_29 <= _GEN_2170;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_30 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_30 <= _GEN_2171;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_31 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_31 <= _GEN_2172;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_32 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_32 <= _GEN_2173;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_33 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_33 <= _GEN_2174;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_34 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_34 <= _GEN_2175;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_35 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_35 <= _GEN_2176;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_36 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_36 <= _GEN_2177;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_37 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_37 <= _GEN_2178;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_38 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_38 <= _GEN_2179;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_39 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_39 <= _GEN_2180;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_40 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_40 <= _GEN_2181;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_41 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_41 <= _GEN_2182;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_42 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_42 <= _GEN_2183;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_43 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_43 <= _GEN_2184;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_44 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_44 <= _GEN_2185;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_45 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_45 <= _GEN_2186;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_46 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_46 <= _GEN_2187;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_47 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_47 <= _GEN_2188;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_48 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_48 <= _GEN_2189;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_49 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_49 <= _GEN_2190;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_50 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_50 <= _GEN_2191;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_51 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_51 <= _GEN_2192;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_52 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_52 <= _GEN_2193;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_53 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_53 <= _GEN_2194;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_54 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_54 <= _GEN_2195;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_55 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_55 <= _GEN_2196;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_56 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_56 <= _GEN_2197;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_57 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_57 <= _GEN_2198;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_58 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_58 <= _GEN_2199;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_59 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_59 <= _GEN_2200;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_60 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_60 <= _GEN_2201;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_61 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_61 <= _GEN_2202;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_62 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_62 <= _GEN_2203;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_63 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_63 <= _GEN_2204;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_64 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_64 <= _GEN_2205;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_65 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_65 <= _GEN_2206;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_66 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_66 <= _GEN_2207;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_67 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_67 <= _GEN_2208;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_68 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_68 <= _GEN_2209;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_69 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_69 <= _GEN_2210;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_70 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_70 <= _GEN_2211;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_71 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_71 <= _GEN_2212;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_72 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_72 <= _GEN_2213;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_73 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_73 <= _GEN_2214;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_74 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_74 <= _GEN_2215;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_75 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_75 <= _GEN_2216;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_76 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_76 <= _GEN_2217;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_77 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_77 <= _GEN_2218;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_78 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_78 <= _GEN_2219;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_79 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_79 <= _GEN_2220;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_80 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_80 <= _GEN_2221;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_81 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_81 <= _GEN_2222;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_82 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_82 <= _GEN_2223;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_83 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_83 <= _GEN_2224;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_84 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_84 <= _GEN_2225;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_85 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_85 <= _GEN_2226;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_86 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_86 <= _GEN_2227;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_87 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_87 <= _GEN_2228;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_88 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_88 <= _GEN_2229;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_89 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_89 <= _GEN_2230;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_90 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_90 <= _GEN_2231;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_91 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_91 <= _GEN_2232;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_92 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_92 <= _GEN_2233;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_93 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_93 <= _GEN_2234;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_94 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_94 <= _GEN_2235;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_95 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_95 <= _GEN_2236;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_96 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_96 <= _GEN_2237;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_97 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_97 <= _GEN_2238;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_98 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_98 <= _GEN_2239;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_99 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_99 <= _GEN_2240;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_100 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_100 <= _GEN_2241;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_101 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_101 <= _GEN_2242;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_102 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_102 <= _GEN_2243;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_103 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_103 <= _GEN_2244;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_104 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_104 <= _GEN_2245;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_105 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_105 <= _GEN_2246;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_106 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_106 <= _GEN_2247;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_107 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_107 <= _GEN_2248;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_108 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_108 <= _GEN_2249;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_109 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_109 <= _GEN_2250;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_110 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_110 <= _GEN_2251;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_111 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_111 <= _GEN_2252;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_112 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_112 <= _GEN_2253;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_113 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_113 <= _GEN_2254;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_114 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_114 <= _GEN_2255;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_115 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_115 <= _GEN_2256;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_116 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_116 <= _GEN_2257;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_117 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_117 <= _GEN_2258;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_118 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_118 <= _GEN_2259;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_119 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_119 <= _GEN_2260;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_120 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_120 <= _GEN_2261;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_121 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_121 <= _GEN_2262;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_122 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_122 <= _GEN_2263;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_123 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_123 <= _GEN_2264;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_124 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_124 <= _GEN_2265;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_125 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_125 <= _GEN_2266;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_126 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_126 <= _GEN_2267;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_127 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_127 <= _GEN_2268;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_128 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_128 <= _GEN_2269;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_129 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_129 <= _GEN_2270;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_130 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_130 <= _GEN_2271;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_131 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_131 <= _GEN_2272;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_132 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_132 <= _GEN_2273;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_133 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_133 <= _GEN_2274;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_134 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_134 <= _GEN_2275;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_135 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_135 <= _GEN_2276;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_136 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_136 <= _GEN_2277;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_137 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_137 <= _GEN_2278;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_138 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_138 <= _GEN_2279;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_139 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_139 <= _GEN_2280;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_140 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_140 <= _GEN_2281;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_141 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_141 <= _GEN_2282;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_142 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_142 <= _GEN_2283;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_143 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_143 <= _GEN_2284;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_144 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_144 <= _GEN_2285;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_145 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_145 <= _GEN_2286;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_146 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_146 <= _GEN_2287;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_147 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_147 <= _GEN_2288;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_148 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_148 <= _GEN_2289;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_149 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_149 <= _GEN_2290;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_150 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_150 <= _GEN_2291;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_151 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_151 <= _GEN_2292;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_152 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_152 <= _GEN_2293;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_153 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_153 <= _GEN_2294;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_154 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_154 <= _GEN_2295;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_155 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_155 <= _GEN_2296;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_156 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_156 <= _GEN_2297;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_157 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_157 <= _GEN_2298;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_158 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_158 <= _GEN_2299;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_159 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_159 <= _GEN_2300;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_160 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_160 <= _GEN_2301;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_161 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_161 <= _GEN_2302;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_162 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_162 <= _GEN_2303;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_163 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_163 <= _GEN_2304;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_164 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_164 <= _GEN_2305;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_165 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_165 <= _GEN_2306;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_166 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_166 <= _GEN_2307;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_167 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_167 <= _GEN_2308;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_168 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_168 <= _GEN_2309;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_169 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_169 <= _GEN_2310;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_170 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_170 <= _GEN_2311;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_171 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_171 <= _GEN_2312;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_172 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_172 <= _GEN_2313;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_173 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_173 <= _GEN_2314;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_174 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_174 <= _GEN_2315;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_175 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_175 <= _GEN_2316;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_176 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_176 <= _GEN_2317;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_177 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_177 <= _GEN_2318;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_178 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_178 <= _GEN_2319;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_179 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_179 <= _GEN_2320;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_180 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_180 <= _GEN_2321;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_181 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_181 <= _GEN_2322;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_182 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_182 <= _GEN_2323;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_183 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_183 <= _GEN_2324;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_184 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_184 <= _GEN_2325;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_185 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_185 <= _GEN_2326;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_186 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_186 <= _GEN_2327;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_187 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_187 <= _GEN_2328;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_188 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_188 <= _GEN_2329;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_189 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_189 <= _GEN_2330;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_190 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_190 <= _GEN_2331;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_191 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_191 <= _GEN_2332;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_192 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_192 <= _GEN_2333;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_193 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_193 <= _GEN_2334;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_194 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_194 <= _GEN_2335;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_195 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_195 <= _GEN_2336;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_196 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_196 <= _GEN_2337;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_197 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_197 <= _GEN_2338;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_198 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_198 <= _GEN_2339;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_199 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_199 <= _GEN_2340;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_200 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_200 <= _GEN_2341;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_201 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_201 <= _GEN_2342;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_202 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_202 <= _GEN_2343;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_203 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_203 <= _GEN_2344;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_204 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_204 <= _GEN_2345;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_205 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_205 <= _GEN_2346;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_206 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_206 <= _GEN_2347;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_207 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_207 <= _GEN_2348;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_208 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_208 <= _GEN_2349;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_209 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_209 <= _GEN_2350;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_210 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_210 <= _GEN_2351;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_211 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_211 <= _GEN_2352;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_212 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_212 <= _GEN_2353;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_213 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_213 <= _GEN_2354;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_214 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_214 <= _GEN_2355;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_215 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_215 <= _GEN_2356;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_216 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_216 <= _GEN_2357;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_217 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_217 <= _GEN_2358;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_218 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_218 <= _GEN_2359;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_219 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_219 <= _GEN_2360;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_220 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_220 <= _GEN_2361;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_221 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_221 <= _GEN_2362;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_222 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_222 <= _GEN_2363;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_223 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_223 <= _GEN_2364;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_224 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_224 <= _GEN_2365;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_225 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_225 <= _GEN_2366;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_226 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_226 <= _GEN_2367;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_227 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_227 <= _GEN_2368;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_228 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_228 <= _GEN_2369;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_229 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_229 <= _GEN_2370;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_230 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_230 <= _GEN_2371;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_231 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_231 <= _GEN_2372;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_232 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_232 <= _GEN_2373;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_233 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_233 <= _GEN_2374;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_234 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_234 <= _GEN_2375;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_235 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_235 <= _GEN_2376;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_236 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_236 <= _GEN_2377;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_237 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_237 <= _GEN_2378;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_238 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_238 <= _GEN_2379;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_239 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_239 <= _GEN_2380;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_240 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_240 <= _GEN_2381;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_241 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_241 <= _GEN_2382;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_242 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_242 <= _GEN_2383;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_243 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_243 <= _GEN_2384;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_244 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_244 <= _GEN_2385;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_245 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_245 <= _GEN_2386;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_246 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_246 <= _GEN_2387;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_247 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_247 <= _GEN_2388;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_248 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_248 <= _GEN_2389;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_249 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_249 <= _GEN_2390;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_250 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_250 <= _GEN_2391;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_251 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_251 <= _GEN_2392;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_252 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_252 <= _GEN_2393;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_253 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_253 <= _GEN_2394;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_254 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_254 <= _GEN_2395;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_255 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_255 <= _GEN_2396;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_256 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_256 <= _GEN_2397;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_257 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_257 <= _GEN_2398;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_258 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_258 <= _GEN_2399;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_259 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_259 <= _GEN_2400;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_260 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_260 <= _GEN_2401;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_261 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_261 <= _GEN_2402;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_262 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_262 <= _GEN_2403;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_263 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_263 <= _GEN_2404;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_264 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_264 <= _GEN_2405;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_265 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_265 <= _GEN_2406;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_266 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_266 <= _GEN_2407;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_267 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_267 <= _GEN_2408;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_268 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_268 <= _GEN_2409;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_269 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_269 <= _GEN_2410;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_270 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_270 <= _GEN_2411;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_271 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_271 <= _GEN_2412;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_272 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_272 <= _GEN_2413;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_273 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_273 <= _GEN_2414;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_274 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_274 <= _GEN_2415;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_275 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_275 <= _GEN_2416;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_276 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_276 <= _GEN_2417;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_277 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_277 <= _GEN_2418;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_278 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_278 <= _GEN_2419;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_279 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_279 <= _GEN_2420;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_280 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_280 <= _GEN_2421;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_281 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_281 <= _GEN_2422;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_282 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_282 <= _GEN_2423;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_283 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_283 <= _GEN_2424;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_284 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_284 <= _GEN_2425;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_285 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_285 <= _GEN_2426;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_286 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_286 <= _GEN_2427;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_287 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_287 <= _GEN_2428;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_288 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_288 <= _GEN_2429;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_289 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_289 <= _GEN_2430;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_290 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_290 <= _GEN_2431;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_291 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_291 <= _GEN_2432;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_292 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_292 <= _GEN_2433;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_293 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_293 <= _GEN_2434;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_294 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_294 <= _GEN_2435;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_295 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_295 <= _GEN_2436;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_296 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_296 <= _GEN_2437;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_297 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_297 <= _GEN_2438;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_298 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_298 <= _GEN_2439;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_299 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_299 <= _GEN_2440;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_300 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_300 <= _GEN_2441;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_301 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_301 <= _GEN_2442;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_302 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_302 <= _GEN_2443;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_303 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_303 <= _GEN_2444;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_304 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_304 <= _GEN_2445;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_305 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_305 <= _GEN_2446;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_306 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_306 <= _GEN_2447;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_307 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_307 <= _GEN_2448;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_308 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_308 <= _GEN_2449;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_309 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_309 <= _GEN_2450;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_310 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_310 <= _GEN_2451;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_311 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_311 <= _GEN_2452;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_312 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_312 <= _GEN_2453;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_313 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_313 <= _GEN_2454;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_314 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_314 <= _GEN_2455;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_315 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_315 <= _GEN_2456;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_316 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_316 <= _GEN_2457;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_317 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_317 <= _GEN_2458;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_318 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_318 <= _GEN_2459;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_319 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_319 <= _GEN_2460;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_320 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_320 <= _GEN_2461;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_321 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_321 <= _GEN_2462;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_322 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_322 <= _GEN_2463;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_323 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_323 <= _GEN_2464;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_324 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_324 <= _GEN_2465;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_325 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_325 <= _GEN_2466;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_326 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_326 <= _GEN_2467;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_327 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_327 <= _GEN_2468;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_328 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_328 <= _GEN_2469;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_329 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_329 <= _GEN_2470;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_330 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_330 <= _GEN_2471;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_331 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_331 <= _GEN_2472;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_332 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_332 <= _GEN_2473;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_333 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_333 <= _GEN_2474;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_334 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_334 <= _GEN_2475;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_335 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_335 <= _GEN_2476;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_336 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_336 <= _GEN_2477;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_337 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_337 <= _GEN_2478;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_338 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_338 <= _GEN_2479;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_339 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_339 <= _GEN_2480;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_340 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_340 <= _GEN_2481;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_341 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_341 <= _GEN_2482;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_342 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_342 <= _GEN_2483;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_343 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_343 <= _GEN_2484;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_344 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_344 <= _GEN_2485;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_345 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_345 <= _GEN_2486;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_346 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_346 <= _GEN_2487;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_347 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_347 <= _GEN_2488;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_348 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_348 <= _GEN_2489;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_349 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_349 <= _GEN_2490;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_350 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_350 <= _GEN_2491;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_351 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_351 <= _GEN_2492;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_352 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_352 <= _GEN_2493;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_353 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_353 <= _GEN_2494;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_354 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_354 <= _GEN_2495;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_355 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_355 <= _GEN_2496;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_356 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_356 <= _GEN_2497;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_357 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_357 <= _GEN_2498;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_358 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_358 <= _GEN_2499;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_359 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_359 <= _GEN_2500;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_360 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_360 <= _GEN_2501;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_361 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_361 <= _GEN_2502;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_362 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_362 <= _GEN_2503;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_363 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_363 <= _GEN_2504;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_364 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_364 <= _GEN_2505;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_365 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_365 <= _GEN_2506;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_366 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_366 <= _GEN_2507;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_367 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_367 <= _GEN_2508;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_368 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_368 <= _GEN_2509;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_369 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_369 <= _GEN_2510;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_370 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_370 <= _GEN_2511;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_371 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_371 <= _GEN_2512;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_372 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_372 <= _GEN_2513;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_373 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_373 <= _GEN_2514;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_374 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_374 <= _GEN_2515;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_375 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_375 <= _GEN_2516;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_376 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_376 <= _GEN_2517;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_377 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_377 <= _GEN_2518;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_378 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_378 <= _GEN_2519;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_379 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_379 <= _GEN_2520;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_380 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_380 <= _GEN_2521;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_381 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_381 <= _GEN_2522;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_382 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_382 <= _GEN_2523;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_383 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_383 <= _GEN_2524;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_384 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_384 <= _GEN_2525;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_385 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_385 <= _GEN_2526;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_386 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_386 <= _GEN_2527;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_387 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_387 <= _GEN_2528;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_388 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_388 <= _GEN_2529;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_389 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_389 <= _GEN_2530;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_390 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_390 <= _GEN_2531;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_391 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_391 <= _GEN_2532;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_392 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_392 <= _GEN_2533;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_393 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_393 <= _GEN_2534;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_394 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_394 <= _GEN_2535;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_395 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_395 <= _GEN_2536;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_396 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_396 <= _GEN_2537;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_397 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_397 <= _GEN_2538;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_398 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_398 <= _GEN_2539;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_399 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_399 <= _GEN_2540;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_400 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_400 <= _GEN_2541;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_401 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_401 <= _GEN_2542;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_402 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_402 <= _GEN_2543;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_403 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_403 <= _GEN_2544;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_404 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_404 <= _GEN_2545;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_405 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_405 <= _GEN_2546;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_406 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_406 <= _GEN_2547;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_407 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_407 <= _GEN_2548;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_408 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_408 <= _GEN_2549;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_409 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_409 <= _GEN_2550;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_410 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_410 <= _GEN_2551;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_411 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_411 <= _GEN_2552;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_412 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_412 <= _GEN_2553;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_413 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_413 <= _GEN_2554;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_414 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_414 <= _GEN_2555;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_415 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_415 <= _GEN_2556;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_416 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_416 <= _GEN_2557;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_417 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_417 <= _GEN_2558;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_418 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_418 <= _GEN_2559;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_419 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_419 <= _GEN_2560;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_420 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_420 <= _GEN_2561;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_421 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_421 <= _GEN_2562;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_422 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_422 <= _GEN_2563;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_423 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_423 <= _GEN_2564;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_424 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_424 <= _GEN_2565;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_425 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_425 <= _GEN_2566;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_426 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_426 <= _GEN_2567;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_427 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_427 <= _GEN_2568;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_428 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_428 <= _GEN_2569;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_429 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_429 <= _GEN_2570;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_430 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_430 <= _GEN_2571;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_431 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_431 <= _GEN_2572;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_432 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_432 <= _GEN_2573;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_433 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_433 <= _GEN_2574;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_434 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_434 <= _GEN_2575;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_435 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_435 <= _GEN_2576;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_436 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_436 <= _GEN_2577;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_437 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_437 <= _GEN_2578;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_438 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_438 <= _GEN_2579;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_439 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_439 <= _GEN_2580;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_440 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_440 <= _GEN_2581;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_441 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_441 <= _GEN_2582;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_442 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_442 <= _GEN_2583;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_443 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_443 <= _GEN_2584;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_444 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_444 <= _GEN_2585;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_445 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_445 <= _GEN_2586;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_446 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_446 <= _GEN_2587;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_447 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_447 <= _GEN_2588;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_448 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_448 <= _GEN_2589;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_449 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_449 <= _GEN_2590;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_450 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_450 <= _GEN_2591;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_451 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_451 <= _GEN_2592;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_452 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_452 <= _GEN_2593;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_453 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_453 <= _GEN_2594;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_454 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_454 <= _GEN_2595;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_455 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_455 <= _GEN_2596;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_456 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_456 <= _GEN_2597;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_457 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_457 <= _GEN_2598;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_458 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_458 <= _GEN_2599;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_459 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_459 <= _GEN_2600;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_460 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_460 <= _GEN_2601;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_461 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_461 <= _GEN_2602;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_462 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_462 <= _GEN_2603;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_463 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_463 <= _GEN_2604;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_464 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_464 <= _GEN_2605;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_465 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_465 <= _GEN_2606;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_466 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_466 <= _GEN_2607;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_467 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_467 <= _GEN_2608;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_468 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_468 <= _GEN_2609;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_469 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_469 <= _GEN_2610;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_470 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_470 <= _GEN_2611;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_471 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_471 <= _GEN_2612;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_472 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_472 <= _GEN_2613;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_473 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_473 <= _GEN_2614;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_474 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_474 <= _GEN_2615;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_475 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_475 <= _GEN_2616;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_476 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_476 <= _GEN_2617;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_477 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_477 <= _GEN_2618;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_478 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_478 <= _GEN_2619;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_479 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_479 <= _GEN_2620;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_480 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_480 <= _GEN_2621;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_481 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_481 <= _GEN_2622;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_482 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_482 <= _GEN_2623;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_483 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_483 <= _GEN_2624;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_484 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_484 <= _GEN_2625;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_485 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_485 <= _GEN_2626;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_486 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_486 <= _GEN_2627;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_487 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_487 <= _GEN_2628;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_488 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_488 <= _GEN_2629;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_489 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_489 <= _GEN_2630;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_490 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_490 <= _GEN_2631;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_491 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_491 <= _GEN_2632;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_492 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_492 <= _GEN_2633;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_493 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_493 <= _GEN_2634;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_494 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_494 <= _GEN_2635;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_495 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_495 <= _GEN_2636;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_496 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_496 <= _GEN_2637;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_497 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_497 <= _GEN_2638;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_498 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_498 <= _GEN_2639;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_499 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_499 <= _GEN_2640;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_500 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_500 <= _GEN_2641;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_501 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_501 <= _GEN_2642;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_502 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_502 <= _GEN_2643;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_503 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_503 <= _GEN_2644;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_504 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_504 <= _GEN_2645;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_505 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_505 <= _GEN_2646;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_506 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_506 <= _GEN_2647;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_507 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_507 <= _GEN_2648;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_508 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_508 <= _GEN_2649;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_509 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_509 <= _GEN_2650;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_510 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_510 <= _GEN_2651;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_511 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_511 <= _GEN_2652;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_512 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_512 <= _GEN_2653;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_513 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_513 <= _GEN_2654;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_514 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_514 <= _GEN_2655;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_515 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_515 <= _GEN_2656;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_516 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_516 <= _GEN_2657;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_517 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_517 <= _GEN_2658;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_518 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_518 <= _GEN_2659;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_519 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_519 <= _GEN_2660;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_520 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_520 <= _GEN_2661;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_521 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_521 <= _GEN_2662;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_522 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_522 <= _GEN_2663;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_523 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_523 <= _GEN_2664;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_524 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_524 <= _GEN_2665;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_525 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_525 <= _GEN_2666;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_526 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_526 <= _GEN_2667;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_527 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_527 <= _GEN_2668;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_528 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_528 <= _GEN_2669;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_529 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_529 <= _GEN_2670;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_530 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_530 <= _GEN_2671;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_531 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_531 <= _GEN_2672;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_532 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_532 <= _GEN_2673;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_533 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_533 <= _GEN_2674;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_534 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_534 <= _GEN_2675;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_535 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_535 <= _GEN_2676;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_536 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_536 <= _GEN_2677;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_537 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_537 <= _GEN_2678;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_538 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_538 <= _GEN_2679;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_539 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_539 <= _GEN_2680;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_540 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_540 <= _GEN_2681;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_541 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_541 <= _GEN_2682;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_542 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_542 <= _GEN_2683;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_543 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_543 <= _GEN_2684;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_544 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_544 <= _GEN_2685;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_545 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_545 <= _GEN_2686;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_546 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_546 <= _GEN_2687;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_547 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_547 <= _GEN_2688;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_548 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_548 <= _GEN_2689;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_549 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_549 <= _GEN_2690;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_550 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_550 <= _GEN_2691;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_551 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_551 <= _GEN_2692;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_552 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_552 <= _GEN_2693;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_553 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_553 <= _GEN_2694;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_554 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_554 <= _GEN_2695;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_555 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_555 <= _GEN_2696;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_556 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_556 <= _GEN_2697;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_557 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_557 <= _GEN_2698;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_558 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_558 <= _GEN_2699;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_559 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_559 <= _GEN_2700;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_560 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_560 <= _GEN_2701;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_561 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_561 <= _GEN_2702;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_562 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_562 <= _GEN_2703;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_563 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_563 <= _GEN_2704;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_564 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_564 <= _GEN_2705;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_565 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_565 <= _GEN_2706;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_566 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_566 <= _GEN_2707;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_567 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_567 <= _GEN_2708;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_568 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_568 <= _GEN_2709;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_569 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_569 <= _GEN_2710;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_570 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_570 <= _GEN_2711;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_571 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_571 <= _GEN_2712;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_572 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_572 <= _GEN_2713;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_573 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_573 <= _GEN_2714;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_574 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_574 <= _GEN_2715;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_575 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_575 <= _GEN_2716;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_576 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_576 <= _GEN_2717;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_577 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_577 <= _GEN_2718;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_578 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_578 <= _GEN_2719;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_579 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_579 <= _GEN_2720;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_580 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_580 <= _GEN_2721;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_581 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_581 <= _GEN_2722;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_582 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_582 <= _GEN_2723;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_583 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_583 <= _GEN_2724;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_584 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_584 <= _GEN_2725;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_585 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_585 <= _GEN_2726;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_586 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_586 <= _GEN_2727;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_587 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_587 <= _GEN_2728;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_588 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_588 <= _GEN_2729;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_589 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_589 <= _GEN_2730;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_590 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_590 <= _GEN_2731;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_591 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_591 <= _GEN_2732;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_592 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_592 <= _GEN_2733;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_593 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_593 <= _GEN_2734;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_594 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_594 <= _GEN_2735;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_595 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_595 <= _GEN_2736;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_596 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_596 <= _GEN_2737;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_597 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_597 <= _GEN_2738;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_598 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_598 <= _GEN_2739;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_599 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_599 <= _GEN_2740;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_600 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_600 <= _GEN_2741;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_601 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_601 <= _GEN_2742;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_602 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_602 <= _GEN_2743;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_603 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_603 <= _GEN_2744;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_604 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_604 <= _GEN_2745;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_605 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_605 <= _GEN_2746;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_606 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_606 <= _GEN_2747;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_607 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_607 <= _GEN_2748;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_608 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_608 <= _GEN_2749;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_609 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_609 <= _GEN_2750;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_610 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_610 <= _GEN_2751;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_611 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_611 <= _GEN_2752;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_612 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_612 <= _GEN_2753;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_613 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_613 <= _GEN_2754;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_614 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_614 <= _GEN_2755;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_615 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_615 <= _GEN_2756;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_616 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_616 <= _GEN_2757;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_617 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_617 <= _GEN_2758;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_618 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_618 <= _GEN_2759;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_619 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_619 <= _GEN_2760;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_620 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_620 <= _GEN_2761;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_621 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_621 <= _GEN_2762;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_622 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_622 <= _GEN_2763;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_623 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_623 <= _GEN_2764;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_624 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_624 <= _GEN_2765;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_625 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_625 <= _GEN_2766;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_626 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_626 <= _GEN_2767;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_627 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_627 <= _GEN_2768;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_628 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_628 <= _GEN_2769;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_629 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_629 <= _GEN_2770;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_630 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_630 <= _GEN_2771;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_631 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_631 <= _GEN_2772;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_632 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_632 <= _GEN_2773;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_633 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_633 <= _GEN_2774;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_634 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_634 <= _GEN_2775;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_635 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_635 <= _GEN_2776;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_636 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_636 <= _GEN_2777;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_637 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_637 <= _GEN_2778;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_638 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_638 <= _GEN_2779;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_639 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_639 <= _GEN_2780;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_640 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_640 <= _GEN_2781;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_641 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_641 <= _GEN_2782;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_642 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_642 <= _GEN_2783;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_643 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_643 <= _GEN_2784;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_644 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_644 <= _GEN_2785;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_645 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_645 <= _GEN_2786;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_646 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_646 <= _GEN_2787;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_647 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_647 <= _GEN_2788;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_648 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_648 <= _GEN_2789;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_649 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_649 <= _GEN_2790;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_650 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_650 <= _GEN_2791;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_651 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_651 <= _GEN_2792;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_652 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_652 <= _GEN_2793;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_653 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_653 <= _GEN_2794;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_654 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_654 <= _GEN_2795;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_655 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_655 <= _GEN_2796;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_656 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_656 <= _GEN_2797;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_657 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_657 <= _GEN_2798;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_658 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_658 <= _GEN_2799;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_659 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_659 <= _GEN_2800;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_660 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_660 <= _GEN_2801;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_661 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_661 <= _GEN_2802;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_662 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_662 <= _GEN_2803;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_663 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_663 <= _GEN_2804;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_664 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_664 <= _GEN_2805;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_665 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_665 <= _GEN_2806;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_666 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_666 <= _GEN_2807;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_667 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_667 <= _GEN_2808;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_668 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_668 <= _GEN_2809;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_669 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_669 <= _GEN_2810;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_670 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_670 <= _GEN_2811;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_671 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_671 <= _GEN_2812;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_672 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_672 <= _GEN_2813;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_673 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_673 <= _GEN_2814;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_674 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_674 <= _GEN_2815;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_675 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_675 <= _GEN_2816;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_676 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_676 <= _GEN_2817;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_677 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_677 <= _GEN_2818;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_678 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_678 <= _GEN_2819;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_679 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_679 <= _GEN_2820;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_680 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_680 <= _GEN_2821;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_681 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_681 <= _GEN_2822;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_682 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_682 <= _GEN_2823;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_683 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_683 <= _GEN_2824;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_684 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_684 <= _GEN_2825;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_685 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_685 <= _GEN_2826;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_686 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_686 <= _GEN_2827;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_687 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_687 <= _GEN_2828;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_688 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_688 <= _GEN_2829;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_689 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_689 <= _GEN_2830;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_690 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_690 <= _GEN_2831;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_691 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_691 <= _GEN_2832;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_692 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_692 <= _GEN_2833;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_693 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_693 <= _GEN_2834;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_694 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_694 <= _GEN_2835;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_695 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_695 <= _GEN_2836;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_696 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_696 <= _GEN_2837;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_697 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_697 <= _GEN_2838;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_698 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_698 <= _GEN_2839;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_699 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_699 <= _GEN_2840;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_700 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_700 <= _GEN_2841;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_701 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_701 <= _GEN_2842;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_702 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_702 <= _GEN_2843;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_703 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_703 <= _GEN_2844;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_704 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_704 <= _GEN_2845;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_705 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_705 <= _GEN_2846;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_706 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_706 <= _GEN_2847;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_707 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_707 <= _GEN_2848;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_708 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_708 <= _GEN_2849;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_709 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_709 <= _GEN_2850;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_710 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_710 <= _GEN_2851;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_711 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_711 <= _GEN_2852;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_712 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_712 <= _GEN_2853;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_713 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_713 <= _GEN_2854;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_714 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_714 <= _GEN_2855;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_715 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_715 <= _GEN_2856;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_716 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_716 <= _GEN_2857;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_717 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_717 <= _GEN_2858;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_718 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_718 <= _GEN_2859;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_719 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_719 <= _GEN_2860;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_720 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_720 <= _GEN_2861;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_721 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_721 <= _GEN_2862;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_722 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_722 <= _GEN_2863;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_723 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_723 <= _GEN_2864;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_724 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_724 <= _GEN_2865;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_725 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_725 <= _GEN_2866;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_726 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_726 <= _GEN_2867;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_727 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_727 <= _GEN_2868;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_728 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_728 <= _GEN_2869;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_729 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_729 <= _GEN_2870;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_730 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_730 <= _GEN_2871;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_731 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_731 <= _GEN_2872;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_732 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_732 <= _GEN_2873;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_733 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_733 <= _GEN_2874;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_734 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_734 <= _GEN_2875;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_735 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_735 <= _GEN_2876;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_736 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_736 <= _GEN_2877;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_737 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_737 <= _GEN_2878;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_738 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_738 <= _GEN_2879;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_739 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_739 <= _GEN_2880;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_740 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_740 <= _GEN_2881;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_741 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_741 <= _GEN_2882;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_742 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_742 <= _GEN_2883;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_743 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_743 <= _GEN_2884;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_744 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_744 <= _GEN_2885;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_745 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_745 <= _GEN_2886;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_746 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_746 <= _GEN_2887;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_747 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_747 <= _GEN_2888;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_748 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_748 <= _GEN_2889;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_749 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_749 <= _GEN_2890;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_750 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_750 <= _GEN_2891;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_751 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_751 <= _GEN_2892;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_752 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_752 <= _GEN_2893;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_753 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_753 <= _GEN_2894;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_754 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_754 <= _GEN_2895;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_755 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_755 <= _GEN_2896;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_756 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_756 <= _GEN_2897;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_757 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_757 <= _GEN_2898;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_758 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_758 <= _GEN_2899;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_759 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_759 <= _GEN_2900;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_760 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_760 <= _GEN_2901;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_761 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_761 <= _GEN_2902;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_762 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_762 <= _GEN_2903;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_763 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_763 <= _GEN_2904;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_764 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_764 <= _GEN_2905;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_765 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_765 <= _GEN_2906;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_766 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_766 <= _GEN_2907;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_767 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_767 <= _GEN_2908;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_768 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_768 <= _GEN_2909;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_769 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_769 <= _GEN_2910;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_770 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_770 <= _GEN_2911;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_771 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_771 <= _GEN_2912;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_772 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_772 <= _GEN_2913;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_773 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_773 <= _GEN_2914;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_774 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_774 <= _GEN_2915;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_775 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_775 <= _GEN_2916;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_776 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_776 <= _GEN_2917;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_777 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_777 <= _GEN_2918;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_778 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_778 <= _GEN_2919;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_779 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_779 <= _GEN_2920;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_780 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_780 <= _GEN_2921;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_781 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_781 <= _GEN_2922;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_782 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_782 <= _GEN_2923;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_783 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_783 <= _GEN_2924;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_784 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_784 <= _GEN_2925;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_785 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_785 <= _GEN_2926;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_786 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_786 <= _GEN_2927;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_787 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_787 <= _GEN_2928;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_788 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_788 <= _GEN_2929;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_789 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_789 <= _GEN_2930;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_790 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_790 <= _GEN_2931;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_791 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_791 <= _GEN_2932;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_792 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_792 <= _GEN_2933;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_793 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_793 <= _GEN_2934;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_794 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_794 <= _GEN_2935;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_795 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_795 <= _GEN_2936;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_796 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_796 <= _GEN_2937;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_797 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_797 <= _GEN_2938;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_798 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_798 <= _GEN_2939;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_799 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_799 <= _GEN_2940;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_800 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_800 <= _GEN_2941;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_801 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_801 <= _GEN_2942;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_802 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_802 <= _GEN_2943;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_803 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_803 <= _GEN_2944;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_804 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_804 <= _GEN_2945;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_805 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_805 <= _GEN_2946;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_806 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_806 <= _GEN_2947;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_807 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_807 <= _GEN_2948;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_808 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_808 <= _GEN_2949;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_809 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_809 <= _GEN_2950;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_810 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_810 <= _GEN_2951;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_811 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_811 <= _GEN_2952;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_812 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_812 <= _GEN_2953;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_813 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_813 <= _GEN_2954;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_814 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_814 <= _GEN_2955;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_815 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_815 <= _GEN_2956;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_816 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_816 <= _GEN_2957;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_817 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_817 <= _GEN_2958;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_818 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_818 <= _GEN_2959;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_819 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_819 <= _GEN_2960;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_820 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_820 <= _GEN_2961;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_821 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_821 <= _GEN_2962;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_822 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_822 <= _GEN_2963;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_823 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_823 <= _GEN_2964;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_824 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_824 <= _GEN_2965;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_825 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_825 <= _GEN_2966;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_826 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_826 <= _GEN_2967;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_827 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_827 <= _GEN_2968;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_828 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_828 <= _GEN_2969;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_829 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_829 <= _GEN_2970;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_830 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_830 <= _GEN_2971;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_831 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_831 <= _GEN_2972;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_832 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_832 <= _GEN_2973;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_833 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_833 <= _GEN_2974;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_834 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_834 <= _GEN_2975;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_835 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_835 <= _GEN_2976;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_836 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_836 <= _GEN_2977;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_837 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_837 <= _GEN_2978;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_838 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_838 <= _GEN_2979;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_839 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_839 <= _GEN_2980;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_840 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_840 <= _GEN_2981;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_841 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_841 <= _GEN_2982;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_842 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_842 <= _GEN_2983;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_843 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_843 <= _GEN_2984;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_844 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_844 <= _GEN_2985;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_845 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_845 <= _GEN_2986;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_846 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_846 <= _GEN_2987;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_847 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_847 <= _GEN_2988;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_848 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_848 <= _GEN_2989;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_849 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_849 <= _GEN_2990;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_850 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_850 <= _GEN_2991;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_851 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_851 <= _GEN_2992;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_852 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_852 <= _GEN_2993;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_853 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_853 <= _GEN_2994;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_854 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_854 <= _GEN_2995;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_855 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_855 <= _GEN_2996;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_856 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_856 <= _GEN_2997;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_857 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_857 <= _GEN_2998;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_858 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_858 <= _GEN_2999;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_859 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_859 <= _GEN_3000;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_860 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_860 <= _GEN_3001;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_861 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_861 <= _GEN_3002;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_862 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_862 <= _GEN_3003;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_863 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_863 <= _GEN_3004;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_864 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_864 <= _GEN_3005;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_865 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_865 <= _GEN_3006;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_866 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_866 <= _GEN_3007;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_867 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_867 <= _GEN_3008;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_868 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_868 <= _GEN_3009;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_869 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_869 <= _GEN_3010;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_870 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_870 <= _GEN_3011;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_871 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_871 <= _GEN_3012;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_872 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_872 <= _GEN_3013;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_873 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_873 <= _GEN_3014;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_874 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_874 <= _GEN_3015;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_875 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_875 <= _GEN_3016;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_876 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_876 <= _GEN_3017;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_877 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_877 <= _GEN_3018;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_878 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_878 <= _GEN_3019;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_879 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_879 <= _GEN_3020;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_880 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_880 <= _GEN_3021;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_881 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_881 <= _GEN_3022;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_882 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_882 <= _GEN_3023;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_883 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_883 <= _GEN_3024;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_884 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_884 <= _GEN_3025;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_885 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_885 <= _GEN_3026;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_886 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_886 <= _GEN_3027;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_887 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_887 <= _GEN_3028;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_888 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_888 <= _GEN_3029;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_889 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_889 <= _GEN_3030;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_890 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_890 <= _GEN_3031;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_891 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_891 <= _GEN_3032;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_892 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_892 <= _GEN_3033;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_893 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_893 <= _GEN_3034;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_894 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_894 <= _GEN_3035;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_895 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_895 <= _GEN_3036;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_896 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_896 <= _GEN_3037;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_897 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_897 <= _GEN_3038;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_898 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_898 <= _GEN_3039;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_899 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_899 <= _GEN_3040;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_900 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_900 <= _GEN_3041;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_901 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_901 <= _GEN_3042;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_902 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_902 <= _GEN_3043;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_903 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_903 <= _GEN_3044;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_904 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_904 <= _GEN_3045;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_905 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_905 <= _GEN_3046;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_906 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_906 <= _GEN_3047;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_907 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_907 <= _GEN_3048;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_908 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_908 <= _GEN_3049;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_909 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_909 <= _GEN_3050;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_910 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_910 <= _GEN_3051;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_911 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_911 <= _GEN_3052;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_912 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_912 <= _GEN_3053;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_913 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_913 <= _GEN_3054;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_914 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_914 <= _GEN_3055;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_915 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_915 <= _GEN_3056;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_916 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_916 <= _GEN_3057;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_917 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_917 <= _GEN_3058;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_918 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_918 <= _GEN_3059;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_919 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_919 <= _GEN_3060;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_920 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_920 <= _GEN_3061;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_921 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_921 <= _GEN_3062;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_922 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_922 <= _GEN_3063;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_923 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_923 <= _GEN_3064;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_924 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_924 <= _GEN_3065;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_925 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_925 <= _GEN_3066;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_926 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_926 <= _GEN_3067;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_927 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_927 <= _GEN_3068;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_928 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_928 <= _GEN_3069;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_929 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_929 <= _GEN_3070;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_930 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_930 <= _GEN_3071;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_931 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_931 <= _GEN_3072;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_932 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_932 <= _GEN_3073;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_933 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_933 <= _GEN_3074;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_934 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_934 <= _GEN_3075;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_935 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_935 <= _GEN_3076;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_936 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_936 <= _GEN_3077;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_937 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_937 <= _GEN_3078;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_938 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_938 <= _GEN_3079;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_939 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_939 <= _GEN_3080;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_940 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_940 <= _GEN_3081;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_941 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_941 <= _GEN_3082;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_942 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_942 <= _GEN_3083;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_943 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_943 <= _GEN_3084;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_944 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_944 <= _GEN_3085;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_945 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_945 <= _GEN_3086;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_946 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_946 <= _GEN_3087;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_947 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_947 <= _GEN_3088;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_948 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_948 <= _GEN_3089;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_949 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_949 <= _GEN_3090;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_950 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_950 <= _GEN_3091;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_951 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_951 <= _GEN_3092;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_952 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_952 <= _GEN_3093;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_953 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_953 <= _GEN_3094;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_954 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_954 <= _GEN_3095;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_955 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_955 <= _GEN_3096;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_956 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_956 <= _GEN_3097;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_957 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_957 <= _GEN_3098;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_958 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_958 <= _GEN_3099;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_959 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_959 <= _GEN_3100;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_960 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_960 <= _GEN_3101;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_961 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_961 <= _GEN_3102;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_962 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_962 <= _GEN_3103;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_963 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_963 <= _GEN_3104;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_964 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_964 <= _GEN_3105;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_965 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_965 <= _GEN_3106;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_966 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_966 <= _GEN_3107;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_967 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_967 <= _GEN_3108;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_968 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_968 <= _GEN_3109;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_969 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_969 <= _GEN_3110;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_970 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_970 <= _GEN_3111;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_971 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_971 <= _GEN_3112;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_972 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_972 <= _GEN_3113;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_973 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_973 <= _GEN_3114;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_974 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_974 <= _GEN_3115;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_975 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_975 <= _GEN_3116;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_976 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_976 <= _GEN_3117;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_977 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_977 <= _GEN_3118;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_978 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_978 <= _GEN_3119;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_979 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_979 <= _GEN_3120;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_980 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_980 <= _GEN_3121;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_981 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_981 <= _GEN_3122;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_982 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_982 <= _GEN_3123;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_983 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_983 <= _GEN_3124;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_984 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_984 <= _GEN_3125;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_985 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_985 <= _GEN_3126;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_986 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_986 <= _GEN_3127;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_987 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_987 <= _GEN_3128;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_988 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_988 <= _GEN_3129;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_989 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_989 <= _GEN_3130;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_990 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_990 <= _GEN_3131;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_991 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_991 <= _GEN_3132;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_992 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_992 <= _GEN_3133;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_993 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_993 <= _GEN_3134;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_994 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_994 <= _GEN_3135;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_995 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_995 <= _GEN_3136;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_996 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_996 <= _GEN_3137;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_997 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_997 <= _GEN_3138;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_998 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_998 <= _GEN_3139;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_999 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_999 <= _GEN_3140;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1000 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1000 <= _GEN_3141;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1001 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1001 <= _GEN_3142;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1002 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1002 <= _GEN_3143;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1003 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1003 <= _GEN_3144;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1004 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1004 <= _GEN_3145;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1005 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1005 <= _GEN_3146;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1006 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1006 <= _GEN_3147;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1007 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1007 <= _GEN_3148;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1008 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1008 <= _GEN_3149;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1009 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1009 <= _GEN_3150;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1010 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1010 <= _GEN_3151;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1011 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1011 <= _GEN_3152;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1012 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1012 <= _GEN_3153;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1013 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1013 <= _GEN_3154;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1014 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1014 <= _GEN_3155;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1015 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1015 <= _GEN_3156;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1016 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1016 <= _GEN_3157;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1017 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1017 <= _GEN_3158;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1018 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1018 <= _GEN_3159;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1019 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1019 <= _GEN_3160;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1020 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1020 <= _GEN_3161;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1021 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1021 <= _GEN_3162;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1022 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1022 <= _GEN_3163;
        end
      end
    end
    if (reset) begin // @[cpu.scala 282:24]
      DMemory_1023 <= 32'h0; // @[cpu.scala 282:24]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (!(_bypassAFromMEM_T_3)) begin // @[cpu.scala 432:29]
        if (!(_stall_T)) begin // @[cpu.scala 434:32]
          DMemory_1023 <= _GEN_3164;
        end
      end
    end
    if (reset) begin // @[cpu.scala 283:24]
      IMemory_0 <= 32'h13; // @[cpu.scala 283:24]
    end else if (io_rvfi_rst) begin // @[cpu.scala 299:21]
      IMemory_0 <= io_rvfi_insn_in_0; // @[cpu.scala 309:18]
    end
    if (reset) begin // @[cpu.scala 283:24]
      IMemory_1 <= 32'h13; // @[cpu.scala 283:24]
    end else if (io_rvfi_rst) begin // @[cpu.scala 299:21]
      IMemory_1 <= io_rvfi_insn_in_1; // @[cpu.scala 309:18]
    end
    if (reset) begin // @[cpu.scala 286:49]
      IFIDIR <= 32'h13; // @[cpu.scala 286:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (~stall) begin // @[cpu.scala 353:27]
        if (~takeBranch) begin // @[cpu.scala 354:34]
          IFIDIR <= ControlUnit_io_insn; // @[cpu.scala 357:16]
        end else begin
          IFIDIR <= 32'h13; // @[cpu.scala 361:16]
        end
      end
    end
    if (reset) begin // @[cpu.scala 286:49]
      IDEXIR <= 32'h13; // @[cpu.scala 286:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (~stall) begin // @[cpu.scala 353:27]
        IDEXIR <= IFIDIR; // @[cpu.scala 406:14]
      end else begin
        IDEXIR <= 32'h13; // @[cpu.scala 408:14]
      end
    end
    if (reset) begin // @[cpu.scala 286:49]
      EXMEMIR <= 32'h13; // @[cpu.scala 286:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      EXMEMIR <= IDEXIR; // @[cpu.scala 428:13]
    end
    if (reset) begin // @[cpu.scala 286:49]
      MEMWBIR <= 32'h13; // @[cpu.scala 286:49]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      MEMWBIR <= EXMEMIR; // @[cpu.scala 440:13]
    end
    if (reset) begin // @[cpu.scala 289:22]
      CurPC <= 64'h0; // @[cpu.scala 289:22]
    end else if (!(io_rvfi_rst)) begin // @[cpu.scala 299:21]
      if (~stall) begin // @[cpu.scala 353:27]
        CurPC <= PC; // @[cpu.scala 377:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  PC = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  Regs_0 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  Regs_1 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  Regs_2 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  Regs_3 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  Regs_4 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  Regs_5 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  Regs_6 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  Regs_7 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  Regs_8 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  Regs_9 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  Regs_10 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  Regs_11 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  Regs_12 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  Regs_13 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  Regs_14 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  Regs_15 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  Regs_16 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  Regs_17 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  Regs_18 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  Regs_19 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  Regs_20 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  Regs_21 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  Regs_22 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  Regs_23 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  Regs_24 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  Regs_25 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  Regs_26 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  Regs_27 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  Regs_28 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  Regs_29 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  Regs_30 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  Regs_31 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  IDEXA = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  IDEXB = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  EXMEMB = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  EXMEMALUOut = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  MEMWBValue = _RAND_37[63:0];
  _RAND_38 = {1{`RANDOM}};
  DMemory_0 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  DMemory_1 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  DMemory_2 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  DMemory_3 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  DMemory_4 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  DMemory_5 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  DMemory_6 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  DMemory_7 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  DMemory_8 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  DMemory_9 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  DMemory_10 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  DMemory_11 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  DMemory_12 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  DMemory_13 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  DMemory_14 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  DMemory_15 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  DMemory_16 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  DMemory_17 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  DMemory_18 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  DMemory_19 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  DMemory_20 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  DMemory_21 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  DMemory_22 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  DMemory_23 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  DMemory_24 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  DMemory_25 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  DMemory_26 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  DMemory_27 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  DMemory_28 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  DMemory_29 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  DMemory_30 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  DMemory_31 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  DMemory_32 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  DMemory_33 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  DMemory_34 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  DMemory_35 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  DMemory_36 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  DMemory_37 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  DMemory_38 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  DMemory_39 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  DMemory_40 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  DMemory_41 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  DMemory_42 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  DMemory_43 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  DMemory_44 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  DMemory_45 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  DMemory_46 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  DMemory_47 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  DMemory_48 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  DMemory_49 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  DMemory_50 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  DMemory_51 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  DMemory_52 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  DMemory_53 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  DMemory_54 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  DMemory_55 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  DMemory_56 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  DMemory_57 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  DMemory_58 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  DMemory_59 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  DMemory_60 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  DMemory_61 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  DMemory_62 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  DMemory_63 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  DMemory_64 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  DMemory_65 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  DMemory_66 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  DMemory_67 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  DMemory_68 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  DMemory_69 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  DMemory_70 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  DMemory_71 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  DMemory_72 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  DMemory_73 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  DMemory_74 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  DMemory_75 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  DMemory_76 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  DMemory_77 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  DMemory_78 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  DMemory_79 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  DMemory_80 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  DMemory_81 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  DMemory_82 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  DMemory_83 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  DMemory_84 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  DMemory_85 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  DMemory_86 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  DMemory_87 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  DMemory_88 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  DMemory_89 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  DMemory_90 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  DMemory_91 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  DMemory_92 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  DMemory_93 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  DMemory_94 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  DMemory_95 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  DMemory_96 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  DMemory_97 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  DMemory_98 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  DMemory_99 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  DMemory_100 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  DMemory_101 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  DMemory_102 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  DMemory_103 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  DMemory_104 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  DMemory_105 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  DMemory_106 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  DMemory_107 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  DMemory_108 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  DMemory_109 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  DMemory_110 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  DMemory_111 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  DMemory_112 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  DMemory_113 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  DMemory_114 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  DMemory_115 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  DMemory_116 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  DMemory_117 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  DMemory_118 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  DMemory_119 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  DMemory_120 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  DMemory_121 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  DMemory_122 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  DMemory_123 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  DMemory_124 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  DMemory_125 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  DMemory_126 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  DMemory_127 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  DMemory_128 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  DMemory_129 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  DMemory_130 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  DMemory_131 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  DMemory_132 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  DMemory_133 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  DMemory_134 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  DMemory_135 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  DMemory_136 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  DMemory_137 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  DMemory_138 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  DMemory_139 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  DMemory_140 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  DMemory_141 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  DMemory_142 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  DMemory_143 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  DMemory_144 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  DMemory_145 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  DMemory_146 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  DMemory_147 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  DMemory_148 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  DMemory_149 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  DMemory_150 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  DMemory_151 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  DMemory_152 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  DMemory_153 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  DMemory_154 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  DMemory_155 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  DMemory_156 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  DMemory_157 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  DMemory_158 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  DMemory_159 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  DMemory_160 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  DMemory_161 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  DMemory_162 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  DMemory_163 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  DMemory_164 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  DMemory_165 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  DMemory_166 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  DMemory_167 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  DMemory_168 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  DMemory_169 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  DMemory_170 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  DMemory_171 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  DMemory_172 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  DMemory_173 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  DMemory_174 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  DMemory_175 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  DMemory_176 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  DMemory_177 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  DMemory_178 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  DMemory_179 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  DMemory_180 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  DMemory_181 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  DMemory_182 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  DMemory_183 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  DMemory_184 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  DMemory_185 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  DMemory_186 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  DMemory_187 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  DMemory_188 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  DMemory_189 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  DMemory_190 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  DMemory_191 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  DMemory_192 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  DMemory_193 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  DMemory_194 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  DMemory_195 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  DMemory_196 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  DMemory_197 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  DMemory_198 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  DMemory_199 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  DMemory_200 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  DMemory_201 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  DMemory_202 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  DMemory_203 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  DMemory_204 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  DMemory_205 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  DMemory_206 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  DMemory_207 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  DMemory_208 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  DMemory_209 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  DMemory_210 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  DMemory_211 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  DMemory_212 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  DMemory_213 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  DMemory_214 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  DMemory_215 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  DMemory_216 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  DMemory_217 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  DMemory_218 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  DMemory_219 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  DMemory_220 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  DMemory_221 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  DMemory_222 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  DMemory_223 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  DMemory_224 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  DMemory_225 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  DMemory_226 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  DMemory_227 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  DMemory_228 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  DMemory_229 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  DMemory_230 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  DMemory_231 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  DMemory_232 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  DMemory_233 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  DMemory_234 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  DMemory_235 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  DMemory_236 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  DMemory_237 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  DMemory_238 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  DMemory_239 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  DMemory_240 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  DMemory_241 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  DMemory_242 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  DMemory_243 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  DMemory_244 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  DMemory_245 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  DMemory_246 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  DMemory_247 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  DMemory_248 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  DMemory_249 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  DMemory_250 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  DMemory_251 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  DMemory_252 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  DMemory_253 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  DMemory_254 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  DMemory_255 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  DMemory_256 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  DMemory_257 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  DMemory_258 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  DMemory_259 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  DMemory_260 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  DMemory_261 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  DMemory_262 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  DMemory_263 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  DMemory_264 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  DMemory_265 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  DMemory_266 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  DMemory_267 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  DMemory_268 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  DMemory_269 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  DMemory_270 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  DMemory_271 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  DMemory_272 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  DMemory_273 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  DMemory_274 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  DMemory_275 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  DMemory_276 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  DMemory_277 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  DMemory_278 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  DMemory_279 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  DMemory_280 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  DMemory_281 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  DMemory_282 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  DMemory_283 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  DMemory_284 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  DMemory_285 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  DMemory_286 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  DMemory_287 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  DMemory_288 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  DMemory_289 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  DMemory_290 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  DMemory_291 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  DMemory_292 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  DMemory_293 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  DMemory_294 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  DMemory_295 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  DMemory_296 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  DMemory_297 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  DMemory_298 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  DMemory_299 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  DMemory_300 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  DMemory_301 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  DMemory_302 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  DMemory_303 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  DMemory_304 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  DMemory_305 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  DMemory_306 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  DMemory_307 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  DMemory_308 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  DMemory_309 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  DMemory_310 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  DMemory_311 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  DMemory_312 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  DMemory_313 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  DMemory_314 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  DMemory_315 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  DMemory_316 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  DMemory_317 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  DMemory_318 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  DMemory_319 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  DMemory_320 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  DMemory_321 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  DMemory_322 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  DMemory_323 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  DMemory_324 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  DMemory_325 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  DMemory_326 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  DMemory_327 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  DMemory_328 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  DMemory_329 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  DMemory_330 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  DMemory_331 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  DMemory_332 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  DMemory_333 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  DMemory_334 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  DMemory_335 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  DMemory_336 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  DMemory_337 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  DMemory_338 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  DMemory_339 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  DMemory_340 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  DMemory_341 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  DMemory_342 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  DMemory_343 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  DMemory_344 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  DMemory_345 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  DMemory_346 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  DMemory_347 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  DMemory_348 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  DMemory_349 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  DMemory_350 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  DMemory_351 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  DMemory_352 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  DMemory_353 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  DMemory_354 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  DMemory_355 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  DMemory_356 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  DMemory_357 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  DMemory_358 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  DMemory_359 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  DMemory_360 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  DMemory_361 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  DMemory_362 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  DMemory_363 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  DMemory_364 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  DMemory_365 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  DMemory_366 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  DMemory_367 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  DMemory_368 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  DMemory_369 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  DMemory_370 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  DMemory_371 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  DMemory_372 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  DMemory_373 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  DMemory_374 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  DMemory_375 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  DMemory_376 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  DMemory_377 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  DMemory_378 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  DMemory_379 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  DMemory_380 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  DMemory_381 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  DMemory_382 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  DMemory_383 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  DMemory_384 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  DMemory_385 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  DMemory_386 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  DMemory_387 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  DMemory_388 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  DMemory_389 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  DMemory_390 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  DMemory_391 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  DMemory_392 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  DMemory_393 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  DMemory_394 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  DMemory_395 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  DMemory_396 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  DMemory_397 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  DMemory_398 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  DMemory_399 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  DMemory_400 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  DMemory_401 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  DMemory_402 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  DMemory_403 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  DMemory_404 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  DMemory_405 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  DMemory_406 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  DMemory_407 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  DMemory_408 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  DMemory_409 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  DMemory_410 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  DMemory_411 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  DMemory_412 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  DMemory_413 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  DMemory_414 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  DMemory_415 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  DMemory_416 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  DMemory_417 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  DMemory_418 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  DMemory_419 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  DMemory_420 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  DMemory_421 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  DMemory_422 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  DMemory_423 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  DMemory_424 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  DMemory_425 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  DMemory_426 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  DMemory_427 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  DMemory_428 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  DMemory_429 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  DMemory_430 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  DMemory_431 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  DMemory_432 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  DMemory_433 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  DMemory_434 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  DMemory_435 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  DMemory_436 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  DMemory_437 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  DMemory_438 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  DMemory_439 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  DMemory_440 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  DMemory_441 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  DMemory_442 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  DMemory_443 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  DMemory_444 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  DMemory_445 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  DMemory_446 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  DMemory_447 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  DMemory_448 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  DMemory_449 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  DMemory_450 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  DMemory_451 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  DMemory_452 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  DMemory_453 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  DMemory_454 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  DMemory_455 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  DMemory_456 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  DMemory_457 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  DMemory_458 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  DMemory_459 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  DMemory_460 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  DMemory_461 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  DMemory_462 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  DMemory_463 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  DMemory_464 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  DMemory_465 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  DMemory_466 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  DMemory_467 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  DMemory_468 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  DMemory_469 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  DMemory_470 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  DMemory_471 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  DMemory_472 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  DMemory_473 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  DMemory_474 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  DMemory_475 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  DMemory_476 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  DMemory_477 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  DMemory_478 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  DMemory_479 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  DMemory_480 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  DMemory_481 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  DMemory_482 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  DMemory_483 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  DMemory_484 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  DMemory_485 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  DMemory_486 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  DMemory_487 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  DMemory_488 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  DMemory_489 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  DMemory_490 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  DMemory_491 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  DMemory_492 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  DMemory_493 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  DMemory_494 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  DMemory_495 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  DMemory_496 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  DMemory_497 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  DMemory_498 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  DMemory_499 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  DMemory_500 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  DMemory_501 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  DMemory_502 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  DMemory_503 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  DMemory_504 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  DMemory_505 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  DMemory_506 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  DMemory_507 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  DMemory_508 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  DMemory_509 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  DMemory_510 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  DMemory_511 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  DMemory_512 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  DMemory_513 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  DMemory_514 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  DMemory_515 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  DMemory_516 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  DMemory_517 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  DMemory_518 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  DMemory_519 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  DMemory_520 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  DMemory_521 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  DMemory_522 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  DMemory_523 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  DMemory_524 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  DMemory_525 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  DMemory_526 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  DMemory_527 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  DMemory_528 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  DMemory_529 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  DMemory_530 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  DMemory_531 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  DMemory_532 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  DMemory_533 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  DMemory_534 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  DMemory_535 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  DMemory_536 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  DMemory_537 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  DMemory_538 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  DMemory_539 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  DMemory_540 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  DMemory_541 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  DMemory_542 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  DMemory_543 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  DMemory_544 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  DMemory_545 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  DMemory_546 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  DMemory_547 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  DMemory_548 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  DMemory_549 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  DMemory_550 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  DMemory_551 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  DMemory_552 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  DMemory_553 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  DMemory_554 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  DMemory_555 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  DMemory_556 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  DMemory_557 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  DMemory_558 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  DMemory_559 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  DMemory_560 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  DMemory_561 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  DMemory_562 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  DMemory_563 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  DMemory_564 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  DMemory_565 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  DMemory_566 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  DMemory_567 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  DMemory_568 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  DMemory_569 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  DMemory_570 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  DMemory_571 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  DMemory_572 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  DMemory_573 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  DMemory_574 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  DMemory_575 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  DMemory_576 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  DMemory_577 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  DMemory_578 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  DMemory_579 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  DMemory_580 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  DMemory_581 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  DMemory_582 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  DMemory_583 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  DMemory_584 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  DMemory_585 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  DMemory_586 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  DMemory_587 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  DMemory_588 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  DMemory_589 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  DMemory_590 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  DMemory_591 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  DMemory_592 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  DMemory_593 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  DMemory_594 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  DMemory_595 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  DMemory_596 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  DMemory_597 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  DMemory_598 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  DMemory_599 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  DMemory_600 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  DMemory_601 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  DMemory_602 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  DMemory_603 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  DMemory_604 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  DMemory_605 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  DMemory_606 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  DMemory_607 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  DMemory_608 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  DMemory_609 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  DMemory_610 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  DMemory_611 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  DMemory_612 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  DMemory_613 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  DMemory_614 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  DMemory_615 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  DMemory_616 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  DMemory_617 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  DMemory_618 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  DMemory_619 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  DMemory_620 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  DMemory_621 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  DMemory_622 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  DMemory_623 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  DMemory_624 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  DMemory_625 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  DMemory_626 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  DMemory_627 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  DMemory_628 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  DMemory_629 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  DMemory_630 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  DMemory_631 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  DMemory_632 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  DMemory_633 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  DMemory_634 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  DMemory_635 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  DMemory_636 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  DMemory_637 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  DMemory_638 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  DMemory_639 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  DMemory_640 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  DMemory_641 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  DMemory_642 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  DMemory_643 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  DMemory_644 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  DMemory_645 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  DMemory_646 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  DMemory_647 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  DMemory_648 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  DMemory_649 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  DMemory_650 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  DMemory_651 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  DMemory_652 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  DMemory_653 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  DMemory_654 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  DMemory_655 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  DMemory_656 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  DMemory_657 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  DMemory_658 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  DMemory_659 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  DMemory_660 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  DMemory_661 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  DMemory_662 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  DMemory_663 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  DMemory_664 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  DMemory_665 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  DMemory_666 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  DMemory_667 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  DMemory_668 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  DMemory_669 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  DMemory_670 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  DMemory_671 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  DMemory_672 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  DMemory_673 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  DMemory_674 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  DMemory_675 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  DMemory_676 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  DMemory_677 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  DMemory_678 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  DMemory_679 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  DMemory_680 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  DMemory_681 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  DMemory_682 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  DMemory_683 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  DMemory_684 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  DMemory_685 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  DMemory_686 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  DMemory_687 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  DMemory_688 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  DMemory_689 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  DMemory_690 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  DMemory_691 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  DMemory_692 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  DMemory_693 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  DMemory_694 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  DMemory_695 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  DMemory_696 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  DMemory_697 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  DMemory_698 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  DMemory_699 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  DMemory_700 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  DMemory_701 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  DMemory_702 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  DMemory_703 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  DMemory_704 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  DMemory_705 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  DMemory_706 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  DMemory_707 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  DMemory_708 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  DMemory_709 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  DMemory_710 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  DMemory_711 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  DMemory_712 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  DMemory_713 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  DMemory_714 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  DMemory_715 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  DMemory_716 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  DMemory_717 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  DMemory_718 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  DMemory_719 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  DMemory_720 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  DMemory_721 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  DMemory_722 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  DMemory_723 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  DMemory_724 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  DMemory_725 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  DMemory_726 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  DMemory_727 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  DMemory_728 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  DMemory_729 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  DMemory_730 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  DMemory_731 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  DMemory_732 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  DMemory_733 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  DMemory_734 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  DMemory_735 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  DMemory_736 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  DMemory_737 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  DMemory_738 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  DMemory_739 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  DMemory_740 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  DMemory_741 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  DMemory_742 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  DMemory_743 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  DMemory_744 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  DMemory_745 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  DMemory_746 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  DMemory_747 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  DMemory_748 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  DMemory_749 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  DMemory_750 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  DMemory_751 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  DMemory_752 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  DMemory_753 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  DMemory_754 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  DMemory_755 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  DMemory_756 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  DMemory_757 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  DMemory_758 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  DMemory_759 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  DMemory_760 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  DMemory_761 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  DMemory_762 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  DMemory_763 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  DMemory_764 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  DMemory_765 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  DMemory_766 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  DMemory_767 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  DMemory_768 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  DMemory_769 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  DMemory_770 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  DMemory_771 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  DMemory_772 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  DMemory_773 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  DMemory_774 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  DMemory_775 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  DMemory_776 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  DMemory_777 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  DMemory_778 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  DMemory_779 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  DMemory_780 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  DMemory_781 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  DMemory_782 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  DMemory_783 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  DMemory_784 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  DMemory_785 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  DMemory_786 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  DMemory_787 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  DMemory_788 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  DMemory_789 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  DMemory_790 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  DMemory_791 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  DMemory_792 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  DMemory_793 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  DMemory_794 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  DMemory_795 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  DMemory_796 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  DMemory_797 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  DMemory_798 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  DMemory_799 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  DMemory_800 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  DMemory_801 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  DMemory_802 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  DMemory_803 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  DMemory_804 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  DMemory_805 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  DMemory_806 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  DMemory_807 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  DMemory_808 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  DMemory_809 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  DMemory_810 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  DMemory_811 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  DMemory_812 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  DMemory_813 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  DMemory_814 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  DMemory_815 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  DMemory_816 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  DMemory_817 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  DMemory_818 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  DMemory_819 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  DMemory_820 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  DMemory_821 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  DMemory_822 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  DMemory_823 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  DMemory_824 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  DMemory_825 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  DMemory_826 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  DMemory_827 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  DMemory_828 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  DMemory_829 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  DMemory_830 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  DMemory_831 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  DMemory_832 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  DMemory_833 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  DMemory_834 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  DMemory_835 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  DMemory_836 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  DMemory_837 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  DMemory_838 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  DMemory_839 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  DMemory_840 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  DMemory_841 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  DMemory_842 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  DMemory_843 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  DMemory_844 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  DMemory_845 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  DMemory_846 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  DMemory_847 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  DMemory_848 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  DMemory_849 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  DMemory_850 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  DMemory_851 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  DMemory_852 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  DMemory_853 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  DMemory_854 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  DMemory_855 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  DMemory_856 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  DMemory_857 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  DMemory_858 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  DMemory_859 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  DMemory_860 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  DMemory_861 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  DMemory_862 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  DMemory_863 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  DMemory_864 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  DMemory_865 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  DMemory_866 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  DMemory_867 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  DMemory_868 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  DMemory_869 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  DMemory_870 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  DMemory_871 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  DMemory_872 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  DMemory_873 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  DMemory_874 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  DMemory_875 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  DMemory_876 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  DMemory_877 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  DMemory_878 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  DMemory_879 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  DMemory_880 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  DMemory_881 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  DMemory_882 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  DMemory_883 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  DMemory_884 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  DMemory_885 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  DMemory_886 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  DMemory_887 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  DMemory_888 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  DMemory_889 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  DMemory_890 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  DMemory_891 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  DMemory_892 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  DMemory_893 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  DMemory_894 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  DMemory_895 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  DMemory_896 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  DMemory_897 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  DMemory_898 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  DMemory_899 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  DMemory_900 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  DMemory_901 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  DMemory_902 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  DMemory_903 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  DMemory_904 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  DMemory_905 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  DMemory_906 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  DMemory_907 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  DMemory_908 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  DMemory_909 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  DMemory_910 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  DMemory_911 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  DMemory_912 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  DMemory_913 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  DMemory_914 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  DMemory_915 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  DMemory_916 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  DMemory_917 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  DMemory_918 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  DMemory_919 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  DMemory_920 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  DMemory_921 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  DMemory_922 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  DMemory_923 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  DMemory_924 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  DMemory_925 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  DMemory_926 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  DMemory_927 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  DMemory_928 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  DMemory_929 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  DMemory_930 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  DMemory_931 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  DMemory_932 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  DMemory_933 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  DMemory_934 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  DMemory_935 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  DMemory_936 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  DMemory_937 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  DMemory_938 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  DMemory_939 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  DMemory_940 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  DMemory_941 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  DMemory_942 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  DMemory_943 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  DMemory_944 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  DMemory_945 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  DMemory_946 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  DMemory_947 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  DMemory_948 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  DMemory_949 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  DMemory_950 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  DMemory_951 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  DMemory_952 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  DMemory_953 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  DMemory_954 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  DMemory_955 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  DMemory_956 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  DMemory_957 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  DMemory_958 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  DMemory_959 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  DMemory_960 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  DMemory_961 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  DMemory_962 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  DMemory_963 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  DMemory_964 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  DMemory_965 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  DMemory_966 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  DMemory_967 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  DMemory_968 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  DMemory_969 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  DMemory_970 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  DMemory_971 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  DMemory_972 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  DMemory_973 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  DMemory_974 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  DMemory_975 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  DMemory_976 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  DMemory_977 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  DMemory_978 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  DMemory_979 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  DMemory_980 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  DMemory_981 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  DMemory_982 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  DMemory_983 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  DMemory_984 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  DMemory_985 = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  DMemory_986 = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  DMemory_987 = _RAND_1025[31:0];
  _RAND_1026 = {1{`RANDOM}};
  DMemory_988 = _RAND_1026[31:0];
  _RAND_1027 = {1{`RANDOM}};
  DMemory_989 = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  DMemory_990 = _RAND_1028[31:0];
  _RAND_1029 = {1{`RANDOM}};
  DMemory_991 = _RAND_1029[31:0];
  _RAND_1030 = {1{`RANDOM}};
  DMemory_992 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  DMemory_993 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  DMemory_994 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  DMemory_995 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  DMemory_996 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  DMemory_997 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  DMemory_998 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  DMemory_999 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  DMemory_1000 = _RAND_1038[31:0];
  _RAND_1039 = {1{`RANDOM}};
  DMemory_1001 = _RAND_1039[31:0];
  _RAND_1040 = {1{`RANDOM}};
  DMemory_1002 = _RAND_1040[31:0];
  _RAND_1041 = {1{`RANDOM}};
  DMemory_1003 = _RAND_1041[31:0];
  _RAND_1042 = {1{`RANDOM}};
  DMemory_1004 = _RAND_1042[31:0];
  _RAND_1043 = {1{`RANDOM}};
  DMemory_1005 = _RAND_1043[31:0];
  _RAND_1044 = {1{`RANDOM}};
  DMemory_1006 = _RAND_1044[31:0];
  _RAND_1045 = {1{`RANDOM}};
  DMemory_1007 = _RAND_1045[31:0];
  _RAND_1046 = {1{`RANDOM}};
  DMemory_1008 = _RAND_1046[31:0];
  _RAND_1047 = {1{`RANDOM}};
  DMemory_1009 = _RAND_1047[31:0];
  _RAND_1048 = {1{`RANDOM}};
  DMemory_1010 = _RAND_1048[31:0];
  _RAND_1049 = {1{`RANDOM}};
  DMemory_1011 = _RAND_1049[31:0];
  _RAND_1050 = {1{`RANDOM}};
  DMemory_1012 = _RAND_1050[31:0];
  _RAND_1051 = {1{`RANDOM}};
  DMemory_1013 = _RAND_1051[31:0];
  _RAND_1052 = {1{`RANDOM}};
  DMemory_1014 = _RAND_1052[31:0];
  _RAND_1053 = {1{`RANDOM}};
  DMemory_1015 = _RAND_1053[31:0];
  _RAND_1054 = {1{`RANDOM}};
  DMemory_1016 = _RAND_1054[31:0];
  _RAND_1055 = {1{`RANDOM}};
  DMemory_1017 = _RAND_1055[31:0];
  _RAND_1056 = {1{`RANDOM}};
  DMemory_1018 = _RAND_1056[31:0];
  _RAND_1057 = {1{`RANDOM}};
  DMemory_1019 = _RAND_1057[31:0];
  _RAND_1058 = {1{`RANDOM}};
  DMemory_1020 = _RAND_1058[31:0];
  _RAND_1059 = {1{`RANDOM}};
  DMemory_1021 = _RAND_1059[31:0];
  _RAND_1060 = {1{`RANDOM}};
  DMemory_1022 = _RAND_1060[31:0];
  _RAND_1061 = {1{`RANDOM}};
  DMemory_1023 = _RAND_1061[31:0];
  _RAND_1062 = {1{`RANDOM}};
  IMemory_0 = _RAND_1062[31:0];
  _RAND_1063 = {1{`RANDOM}};
  IMemory_1 = _RAND_1063[31:0];
  _RAND_1064 = {1{`RANDOM}};
  IFIDIR = _RAND_1064[31:0];
  _RAND_1065 = {1{`RANDOM}};
  IDEXIR = _RAND_1065[31:0];
  _RAND_1066 = {1{`RANDOM}};
  EXMEMIR = _RAND_1066[31:0];
  _RAND_1067 = {1{`RANDOM}};
  MEMWBIR = _RAND_1067[31:0];
  _RAND_1068 = {2{`RANDOM}};
  CurPC = _RAND_1068[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module self(
  input         clock,
  input         reset,
  input  [31:0] io_insn_in_0,
  input  [31:0] io_insn_in_1,
  input  [31:0] io_insn_in_2,
  input  [31:0] io_insn_in_3,
  input  [31:0] io_insn_in_4,
  input  [31:0] io_insn_in_5,
  input  [31:0] io_insn_in_6,
  input  [31:0] io_insn_in_7,
  input         io_rst,
  output        io_o
);
  wire  cpu1_clock; // @[cpu.scala 490:20]
  wire  cpu1_reset; // @[cpu.scala 490:20]
  wire  cpu1_io_rvfi_rst; // @[cpu.scala 490:20]
  wire [31:0] cpu1_io_rvfi_insn_in_0; // @[cpu.scala 490:20]
  wire [31:0] cpu1_io_rvfi_insn_in_1; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_0; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_1; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_2; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_3; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_4; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_5; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_6; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_7; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_8; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_9; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_10; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_11; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_12; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_13; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_14; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_15; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_16; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_17; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_18; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_19; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_20; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_21; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_22; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_23; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_24; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_25; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_26; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_27; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_28; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_29; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_30; // @[cpu.scala 490:20]
  wire [63:0] cpu1_io_rvfi_regs_31; // @[cpu.scala 490:20]
  wire  cpu2_clock; // @[cpu.scala 491:20]
  wire  cpu2_reset; // @[cpu.scala 491:20]
  wire  cpu2_io_rvfi_rst; // @[cpu.scala 491:20]
  wire [31:0] cpu2_io_rvfi_insn_in_0; // @[cpu.scala 491:20]
  wire [31:0] cpu2_io_rvfi_insn_in_1; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_0; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_1; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_2; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_3; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_4; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_5; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_6; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_7; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_8; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_9; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_10; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_11; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_12; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_13; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_14; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_15; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_16; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_17; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_18; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_19; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_20; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_21; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_22; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_23; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_24; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_25; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_26; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_27; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_28; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_29; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_30; // @[cpu.scala 491:20]
  wire [63:0] cpu2_io_rvfi_regs_31; // @[cpu.scala 491:20]
  wire  _equalreg_T_15 = cpu1_io_rvfi_regs_15 == cpu2_io_rvfi_regs_15; // @[cpu.scala 505:82]
  wire  _equalreg_T_46 = cpu1_io_rvfi_regs_0 == cpu2_io_rvfi_regs_0 & cpu1_io_rvfi_regs_1 == cpu2_io_rvfi_regs_1 &
    cpu1_io_rvfi_regs_2 == cpu2_io_rvfi_regs_2 & cpu1_io_rvfi_regs_3 == cpu2_io_rvfi_regs_3 & cpu1_io_rvfi_regs_4 ==
    cpu2_io_rvfi_regs_4 & cpu1_io_rvfi_regs_5 == cpu2_io_rvfi_regs_5 & cpu1_io_rvfi_regs_6 == cpu2_io_rvfi_regs_6 &
    cpu1_io_rvfi_regs_7 == cpu2_io_rvfi_regs_7 & cpu1_io_rvfi_regs_8 == cpu2_io_rvfi_regs_8 & cpu1_io_rvfi_regs_9 ==
    cpu2_io_rvfi_regs_9 & cpu1_io_rvfi_regs_10 == cpu2_io_rvfi_regs_10 & cpu1_io_rvfi_regs_11 == cpu2_io_rvfi_regs_11 &
    cpu1_io_rvfi_regs_12 == cpu2_io_rvfi_regs_12 & cpu1_io_rvfi_regs_13 == cpu2_io_rvfi_regs_13 & cpu1_io_rvfi_regs_14
     == cpu2_io_rvfi_regs_14 & _equalreg_T_15; // @[cpu.scala 505:99]
  wire  _equalreg_T_61 = _equalreg_T_46 & cpu1_io_rvfi_regs_16 == cpu2_io_rvfi_regs_16 & cpu1_io_rvfi_regs_17 ==
    cpu2_io_rvfi_regs_17 & cpu1_io_rvfi_regs_18 == cpu2_io_rvfi_regs_18 & cpu1_io_rvfi_regs_19 == cpu2_io_rvfi_regs_19
     & cpu1_io_rvfi_regs_20 == cpu2_io_rvfi_regs_20 & cpu1_io_rvfi_regs_21 == cpu2_io_rvfi_regs_21 &
    cpu1_io_rvfi_regs_22 == cpu2_io_rvfi_regs_22 & cpu1_io_rvfi_regs_23 == cpu2_io_rvfi_regs_23 & cpu1_io_rvfi_regs_24
     == cpu2_io_rvfi_regs_24 & cpu1_io_rvfi_regs_25 == cpu2_io_rvfi_regs_25 & cpu1_io_rvfi_regs_26 ==
    cpu2_io_rvfi_regs_26 & cpu1_io_rvfi_regs_27 == cpu2_io_rvfi_regs_27 & cpu1_io_rvfi_regs_28 == cpu2_io_rvfi_regs_28
     & cpu1_io_rvfi_regs_29 == cpu2_io_rvfi_regs_29 & cpu1_io_rvfi_regs_30 == cpu2_io_rvfi_regs_30; // @[cpu.scala 505:99]
  RISCVCPUv2 cpu1 ( // @[cpu.scala 490:20]
    .clock(cpu1_clock),
    .reset(cpu1_reset),
    .io_rvfi_rst(cpu1_io_rvfi_rst),
    .io_rvfi_insn_in_0(cpu1_io_rvfi_insn_in_0),
    .io_rvfi_insn_in_1(cpu1_io_rvfi_insn_in_1),
    .io_rvfi_regs_0(cpu1_io_rvfi_regs_0),
    .io_rvfi_regs_1(cpu1_io_rvfi_regs_1),
    .io_rvfi_regs_2(cpu1_io_rvfi_regs_2),
    .io_rvfi_regs_3(cpu1_io_rvfi_regs_3),
    .io_rvfi_regs_4(cpu1_io_rvfi_regs_4),
    .io_rvfi_regs_5(cpu1_io_rvfi_regs_5),
    .io_rvfi_regs_6(cpu1_io_rvfi_regs_6),
    .io_rvfi_regs_7(cpu1_io_rvfi_regs_7),
    .io_rvfi_regs_8(cpu1_io_rvfi_regs_8),
    .io_rvfi_regs_9(cpu1_io_rvfi_regs_9),
    .io_rvfi_regs_10(cpu1_io_rvfi_regs_10),
    .io_rvfi_regs_11(cpu1_io_rvfi_regs_11),
    .io_rvfi_regs_12(cpu1_io_rvfi_regs_12),
    .io_rvfi_regs_13(cpu1_io_rvfi_regs_13),
    .io_rvfi_regs_14(cpu1_io_rvfi_regs_14),
    .io_rvfi_regs_15(cpu1_io_rvfi_regs_15),
    .io_rvfi_regs_16(cpu1_io_rvfi_regs_16),
    .io_rvfi_regs_17(cpu1_io_rvfi_regs_17),
    .io_rvfi_regs_18(cpu1_io_rvfi_regs_18),
    .io_rvfi_regs_19(cpu1_io_rvfi_regs_19),
    .io_rvfi_regs_20(cpu1_io_rvfi_regs_20),
    .io_rvfi_regs_21(cpu1_io_rvfi_regs_21),
    .io_rvfi_regs_22(cpu1_io_rvfi_regs_22),
    .io_rvfi_regs_23(cpu1_io_rvfi_regs_23),
    .io_rvfi_regs_24(cpu1_io_rvfi_regs_24),
    .io_rvfi_regs_25(cpu1_io_rvfi_regs_25),
    .io_rvfi_regs_26(cpu1_io_rvfi_regs_26),
    .io_rvfi_regs_27(cpu1_io_rvfi_regs_27),
    .io_rvfi_regs_28(cpu1_io_rvfi_regs_28),
    .io_rvfi_regs_29(cpu1_io_rvfi_regs_29),
    .io_rvfi_regs_30(cpu1_io_rvfi_regs_30),
    .io_rvfi_regs_31(cpu1_io_rvfi_regs_31)
  );
  RISCVCPUv2Bubble cpu2 ( // @[cpu.scala 491:20]
    .clock(cpu2_clock),
    .reset(cpu2_reset),
    .io_rvfi_rst(cpu2_io_rvfi_rst),
    .io_rvfi_insn_in_0(cpu2_io_rvfi_insn_in_0),
    .io_rvfi_insn_in_1(cpu2_io_rvfi_insn_in_1),
    .io_rvfi_regs_0(cpu2_io_rvfi_regs_0),
    .io_rvfi_regs_1(cpu2_io_rvfi_regs_1),
    .io_rvfi_regs_2(cpu2_io_rvfi_regs_2),
    .io_rvfi_regs_3(cpu2_io_rvfi_regs_3),
    .io_rvfi_regs_4(cpu2_io_rvfi_regs_4),
    .io_rvfi_regs_5(cpu2_io_rvfi_regs_5),
    .io_rvfi_regs_6(cpu2_io_rvfi_regs_6),
    .io_rvfi_regs_7(cpu2_io_rvfi_regs_7),
    .io_rvfi_regs_8(cpu2_io_rvfi_regs_8),
    .io_rvfi_regs_9(cpu2_io_rvfi_regs_9),
    .io_rvfi_regs_10(cpu2_io_rvfi_regs_10),
    .io_rvfi_regs_11(cpu2_io_rvfi_regs_11),
    .io_rvfi_regs_12(cpu2_io_rvfi_regs_12),
    .io_rvfi_regs_13(cpu2_io_rvfi_regs_13),
    .io_rvfi_regs_14(cpu2_io_rvfi_regs_14),
    .io_rvfi_regs_15(cpu2_io_rvfi_regs_15),
    .io_rvfi_regs_16(cpu2_io_rvfi_regs_16),
    .io_rvfi_regs_17(cpu2_io_rvfi_regs_17),
    .io_rvfi_regs_18(cpu2_io_rvfi_regs_18),
    .io_rvfi_regs_19(cpu2_io_rvfi_regs_19),
    .io_rvfi_regs_20(cpu2_io_rvfi_regs_20),
    .io_rvfi_regs_21(cpu2_io_rvfi_regs_21),
    .io_rvfi_regs_22(cpu2_io_rvfi_regs_22),
    .io_rvfi_regs_23(cpu2_io_rvfi_regs_23),
    .io_rvfi_regs_24(cpu2_io_rvfi_regs_24),
    .io_rvfi_regs_25(cpu2_io_rvfi_regs_25),
    .io_rvfi_regs_26(cpu2_io_rvfi_regs_26),
    .io_rvfi_regs_27(cpu2_io_rvfi_regs_27),
    .io_rvfi_regs_28(cpu2_io_rvfi_regs_28),
    .io_rvfi_regs_29(cpu2_io_rvfi_regs_29),
    .io_rvfi_regs_30(cpu2_io_rvfi_regs_30),
    .io_rvfi_regs_31(cpu2_io_rvfi_regs_31)
  );
  assign io_o = _equalreg_T_61 & cpu1_io_rvfi_regs_31 == cpu2_io_rvfi_regs_31; // @[cpu.scala 505:99]
  assign cpu1_clock = clock;
  assign cpu1_reset = reset;
  assign cpu1_io_rvfi_rst = io_rst; // @[cpu.scala 503:20]
  assign cpu1_io_rvfi_insn_in_0 = io_insn_in_0; // @[cpu.scala 494:31]
  assign cpu1_io_rvfi_insn_in_1 = io_insn_in_1; // @[cpu.scala 494:31]
  assign cpu2_clock = clock;
  assign cpu2_reset = reset;
  assign cpu2_io_rvfi_rst = io_rst; // @[cpu.scala 504:20]
  assign cpu2_io_rvfi_insn_in_0 = io_insn_in_0; // @[cpu.scala 495:31]
  assign cpu2_io_rvfi_insn_in_1 = io_insn_in_1; // @[cpu.scala 495:31]
endmodule
