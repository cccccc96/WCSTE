module CAMLine(
  input          clock,
  input          io_we,
  input          io_wi,
  input  [255:0] io_key,
  input  [255:0] io_din,
  output         io_hit
);
`ifdef RANDOMIZE_REG_INIT
  reg [255:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  write = io_we & io_wi; // @[cam.scala 58:18]
  reg [255:0] camCells; // @[cam.scala 59:21]
  assign io_hit = camCells == io_key; // @[cam.scala 65:23]
  always @(posedge clock) begin
    if (write) begin // @[cam.scala 61:14]
      camCells <= io_din; // @[cam.scala 62:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  camCells = _RAND_0[255:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CAM_m_n(
  input          clock,
  input          reset,
  input          io_we,
  input  [255:0] io_key,
  input  [255:0] io_din,
  input  [255:0] io_waddr,
  output         io_hit
);
  wire  CAMLine_clock; // @[cam.scala 81:36]
  wire  CAMLine_io_we; // @[cam.scala 81:36]
  wire  CAMLine_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_io_din; // @[cam.scala 81:36]
  wire  CAMLine_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_1_clock; // @[cam.scala 81:36]
  wire  CAMLine_1_io_we; // @[cam.scala 81:36]
  wire  CAMLine_1_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_1_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_1_io_din; // @[cam.scala 81:36]
  wire  CAMLine_1_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_2_clock; // @[cam.scala 81:36]
  wire  CAMLine_2_io_we; // @[cam.scala 81:36]
  wire  CAMLine_2_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_2_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_2_io_din; // @[cam.scala 81:36]
  wire  CAMLine_2_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_3_clock; // @[cam.scala 81:36]
  wire  CAMLine_3_io_we; // @[cam.scala 81:36]
  wire  CAMLine_3_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_3_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_3_io_din; // @[cam.scala 81:36]
  wire  CAMLine_3_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_4_clock; // @[cam.scala 81:36]
  wire  CAMLine_4_io_we; // @[cam.scala 81:36]
  wire  CAMLine_4_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_4_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_4_io_din; // @[cam.scala 81:36]
  wire  CAMLine_4_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_5_clock; // @[cam.scala 81:36]
  wire  CAMLine_5_io_we; // @[cam.scala 81:36]
  wire  CAMLine_5_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_5_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_5_io_din; // @[cam.scala 81:36]
  wire  CAMLine_5_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_6_clock; // @[cam.scala 81:36]
  wire  CAMLine_6_io_we; // @[cam.scala 81:36]
  wire  CAMLine_6_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_6_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_6_io_din; // @[cam.scala 81:36]
  wire  CAMLine_6_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_7_clock; // @[cam.scala 81:36]
  wire  CAMLine_7_io_we; // @[cam.scala 81:36]
  wire  CAMLine_7_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_7_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_7_io_din; // @[cam.scala 81:36]
  wire  CAMLine_7_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_8_clock; // @[cam.scala 81:36]
  wire  CAMLine_8_io_we; // @[cam.scala 81:36]
  wire  CAMLine_8_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_8_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_8_io_din; // @[cam.scala 81:36]
  wire  CAMLine_8_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_9_clock; // @[cam.scala 81:36]
  wire  CAMLine_9_io_we; // @[cam.scala 81:36]
  wire  CAMLine_9_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_9_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_9_io_din; // @[cam.scala 81:36]
  wire  CAMLine_9_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_10_clock; // @[cam.scala 81:36]
  wire  CAMLine_10_io_we; // @[cam.scala 81:36]
  wire  CAMLine_10_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_10_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_10_io_din; // @[cam.scala 81:36]
  wire  CAMLine_10_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_11_clock; // @[cam.scala 81:36]
  wire  CAMLine_11_io_we; // @[cam.scala 81:36]
  wire  CAMLine_11_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_11_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_11_io_din; // @[cam.scala 81:36]
  wire  CAMLine_11_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_12_clock; // @[cam.scala 81:36]
  wire  CAMLine_12_io_we; // @[cam.scala 81:36]
  wire  CAMLine_12_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_12_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_12_io_din; // @[cam.scala 81:36]
  wire  CAMLine_12_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_13_clock; // @[cam.scala 81:36]
  wire  CAMLine_13_io_we; // @[cam.scala 81:36]
  wire  CAMLine_13_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_13_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_13_io_din; // @[cam.scala 81:36]
  wire  CAMLine_13_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_14_clock; // @[cam.scala 81:36]
  wire  CAMLine_14_io_we; // @[cam.scala 81:36]
  wire  CAMLine_14_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_14_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_14_io_din; // @[cam.scala 81:36]
  wire  CAMLine_14_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_15_clock; // @[cam.scala 81:36]
  wire  CAMLine_15_io_we; // @[cam.scala 81:36]
  wire  CAMLine_15_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_15_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_15_io_din; // @[cam.scala 81:36]
  wire  CAMLine_15_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_16_clock; // @[cam.scala 81:36]
  wire  CAMLine_16_io_we; // @[cam.scala 81:36]
  wire  CAMLine_16_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_16_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_16_io_din; // @[cam.scala 81:36]
  wire  CAMLine_16_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_17_clock; // @[cam.scala 81:36]
  wire  CAMLine_17_io_we; // @[cam.scala 81:36]
  wire  CAMLine_17_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_17_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_17_io_din; // @[cam.scala 81:36]
  wire  CAMLine_17_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_18_clock; // @[cam.scala 81:36]
  wire  CAMLine_18_io_we; // @[cam.scala 81:36]
  wire  CAMLine_18_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_18_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_18_io_din; // @[cam.scala 81:36]
  wire  CAMLine_18_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_19_clock; // @[cam.scala 81:36]
  wire  CAMLine_19_io_we; // @[cam.scala 81:36]
  wire  CAMLine_19_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_19_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_19_io_din; // @[cam.scala 81:36]
  wire  CAMLine_19_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_20_clock; // @[cam.scala 81:36]
  wire  CAMLine_20_io_we; // @[cam.scala 81:36]
  wire  CAMLine_20_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_20_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_20_io_din; // @[cam.scala 81:36]
  wire  CAMLine_20_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_21_clock; // @[cam.scala 81:36]
  wire  CAMLine_21_io_we; // @[cam.scala 81:36]
  wire  CAMLine_21_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_21_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_21_io_din; // @[cam.scala 81:36]
  wire  CAMLine_21_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_22_clock; // @[cam.scala 81:36]
  wire  CAMLine_22_io_we; // @[cam.scala 81:36]
  wire  CAMLine_22_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_22_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_22_io_din; // @[cam.scala 81:36]
  wire  CAMLine_22_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_23_clock; // @[cam.scala 81:36]
  wire  CAMLine_23_io_we; // @[cam.scala 81:36]
  wire  CAMLine_23_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_23_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_23_io_din; // @[cam.scala 81:36]
  wire  CAMLine_23_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_24_clock; // @[cam.scala 81:36]
  wire  CAMLine_24_io_we; // @[cam.scala 81:36]
  wire  CAMLine_24_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_24_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_24_io_din; // @[cam.scala 81:36]
  wire  CAMLine_24_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_25_clock; // @[cam.scala 81:36]
  wire  CAMLine_25_io_we; // @[cam.scala 81:36]
  wire  CAMLine_25_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_25_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_25_io_din; // @[cam.scala 81:36]
  wire  CAMLine_25_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_26_clock; // @[cam.scala 81:36]
  wire  CAMLine_26_io_we; // @[cam.scala 81:36]
  wire  CAMLine_26_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_26_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_26_io_din; // @[cam.scala 81:36]
  wire  CAMLine_26_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_27_clock; // @[cam.scala 81:36]
  wire  CAMLine_27_io_we; // @[cam.scala 81:36]
  wire  CAMLine_27_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_27_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_27_io_din; // @[cam.scala 81:36]
  wire  CAMLine_27_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_28_clock; // @[cam.scala 81:36]
  wire  CAMLine_28_io_we; // @[cam.scala 81:36]
  wire  CAMLine_28_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_28_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_28_io_din; // @[cam.scala 81:36]
  wire  CAMLine_28_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_29_clock; // @[cam.scala 81:36]
  wire  CAMLine_29_io_we; // @[cam.scala 81:36]
  wire  CAMLine_29_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_29_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_29_io_din; // @[cam.scala 81:36]
  wire  CAMLine_29_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_30_clock; // @[cam.scala 81:36]
  wire  CAMLine_30_io_we; // @[cam.scala 81:36]
  wire  CAMLine_30_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_30_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_30_io_din; // @[cam.scala 81:36]
  wire  CAMLine_30_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_31_clock; // @[cam.scala 81:36]
  wire  CAMLine_31_io_we; // @[cam.scala 81:36]
  wire  CAMLine_31_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_31_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_31_io_din; // @[cam.scala 81:36]
  wire  CAMLine_31_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_32_clock; // @[cam.scala 81:36]
  wire  CAMLine_32_io_we; // @[cam.scala 81:36]
  wire  CAMLine_32_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_32_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_32_io_din; // @[cam.scala 81:36]
  wire  CAMLine_32_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_33_clock; // @[cam.scala 81:36]
  wire  CAMLine_33_io_we; // @[cam.scala 81:36]
  wire  CAMLine_33_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_33_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_33_io_din; // @[cam.scala 81:36]
  wire  CAMLine_33_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_34_clock; // @[cam.scala 81:36]
  wire  CAMLine_34_io_we; // @[cam.scala 81:36]
  wire  CAMLine_34_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_34_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_34_io_din; // @[cam.scala 81:36]
  wire  CAMLine_34_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_35_clock; // @[cam.scala 81:36]
  wire  CAMLine_35_io_we; // @[cam.scala 81:36]
  wire  CAMLine_35_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_35_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_35_io_din; // @[cam.scala 81:36]
  wire  CAMLine_35_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_36_clock; // @[cam.scala 81:36]
  wire  CAMLine_36_io_we; // @[cam.scala 81:36]
  wire  CAMLine_36_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_36_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_36_io_din; // @[cam.scala 81:36]
  wire  CAMLine_36_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_37_clock; // @[cam.scala 81:36]
  wire  CAMLine_37_io_we; // @[cam.scala 81:36]
  wire  CAMLine_37_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_37_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_37_io_din; // @[cam.scala 81:36]
  wire  CAMLine_37_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_38_clock; // @[cam.scala 81:36]
  wire  CAMLine_38_io_we; // @[cam.scala 81:36]
  wire  CAMLine_38_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_38_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_38_io_din; // @[cam.scala 81:36]
  wire  CAMLine_38_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_39_clock; // @[cam.scala 81:36]
  wire  CAMLine_39_io_we; // @[cam.scala 81:36]
  wire  CAMLine_39_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_39_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_39_io_din; // @[cam.scala 81:36]
  wire  CAMLine_39_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_40_clock; // @[cam.scala 81:36]
  wire  CAMLine_40_io_we; // @[cam.scala 81:36]
  wire  CAMLine_40_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_40_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_40_io_din; // @[cam.scala 81:36]
  wire  CAMLine_40_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_41_clock; // @[cam.scala 81:36]
  wire  CAMLine_41_io_we; // @[cam.scala 81:36]
  wire  CAMLine_41_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_41_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_41_io_din; // @[cam.scala 81:36]
  wire  CAMLine_41_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_42_clock; // @[cam.scala 81:36]
  wire  CAMLine_42_io_we; // @[cam.scala 81:36]
  wire  CAMLine_42_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_42_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_42_io_din; // @[cam.scala 81:36]
  wire  CAMLine_42_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_43_clock; // @[cam.scala 81:36]
  wire  CAMLine_43_io_we; // @[cam.scala 81:36]
  wire  CAMLine_43_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_43_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_43_io_din; // @[cam.scala 81:36]
  wire  CAMLine_43_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_44_clock; // @[cam.scala 81:36]
  wire  CAMLine_44_io_we; // @[cam.scala 81:36]
  wire  CAMLine_44_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_44_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_44_io_din; // @[cam.scala 81:36]
  wire  CAMLine_44_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_45_clock; // @[cam.scala 81:36]
  wire  CAMLine_45_io_we; // @[cam.scala 81:36]
  wire  CAMLine_45_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_45_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_45_io_din; // @[cam.scala 81:36]
  wire  CAMLine_45_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_46_clock; // @[cam.scala 81:36]
  wire  CAMLine_46_io_we; // @[cam.scala 81:36]
  wire  CAMLine_46_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_46_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_46_io_din; // @[cam.scala 81:36]
  wire  CAMLine_46_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_47_clock; // @[cam.scala 81:36]
  wire  CAMLine_47_io_we; // @[cam.scala 81:36]
  wire  CAMLine_47_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_47_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_47_io_din; // @[cam.scala 81:36]
  wire  CAMLine_47_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_48_clock; // @[cam.scala 81:36]
  wire  CAMLine_48_io_we; // @[cam.scala 81:36]
  wire  CAMLine_48_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_48_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_48_io_din; // @[cam.scala 81:36]
  wire  CAMLine_48_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_49_clock; // @[cam.scala 81:36]
  wire  CAMLine_49_io_we; // @[cam.scala 81:36]
  wire  CAMLine_49_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_49_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_49_io_din; // @[cam.scala 81:36]
  wire  CAMLine_49_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_50_clock; // @[cam.scala 81:36]
  wire  CAMLine_50_io_we; // @[cam.scala 81:36]
  wire  CAMLine_50_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_50_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_50_io_din; // @[cam.scala 81:36]
  wire  CAMLine_50_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_51_clock; // @[cam.scala 81:36]
  wire  CAMLine_51_io_we; // @[cam.scala 81:36]
  wire  CAMLine_51_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_51_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_51_io_din; // @[cam.scala 81:36]
  wire  CAMLine_51_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_52_clock; // @[cam.scala 81:36]
  wire  CAMLine_52_io_we; // @[cam.scala 81:36]
  wire  CAMLine_52_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_52_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_52_io_din; // @[cam.scala 81:36]
  wire  CAMLine_52_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_53_clock; // @[cam.scala 81:36]
  wire  CAMLine_53_io_we; // @[cam.scala 81:36]
  wire  CAMLine_53_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_53_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_53_io_din; // @[cam.scala 81:36]
  wire  CAMLine_53_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_54_clock; // @[cam.scala 81:36]
  wire  CAMLine_54_io_we; // @[cam.scala 81:36]
  wire  CAMLine_54_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_54_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_54_io_din; // @[cam.scala 81:36]
  wire  CAMLine_54_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_55_clock; // @[cam.scala 81:36]
  wire  CAMLine_55_io_we; // @[cam.scala 81:36]
  wire  CAMLine_55_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_55_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_55_io_din; // @[cam.scala 81:36]
  wire  CAMLine_55_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_56_clock; // @[cam.scala 81:36]
  wire  CAMLine_56_io_we; // @[cam.scala 81:36]
  wire  CAMLine_56_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_56_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_56_io_din; // @[cam.scala 81:36]
  wire  CAMLine_56_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_57_clock; // @[cam.scala 81:36]
  wire  CAMLine_57_io_we; // @[cam.scala 81:36]
  wire  CAMLine_57_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_57_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_57_io_din; // @[cam.scala 81:36]
  wire  CAMLine_57_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_58_clock; // @[cam.scala 81:36]
  wire  CAMLine_58_io_we; // @[cam.scala 81:36]
  wire  CAMLine_58_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_58_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_58_io_din; // @[cam.scala 81:36]
  wire  CAMLine_58_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_59_clock; // @[cam.scala 81:36]
  wire  CAMLine_59_io_we; // @[cam.scala 81:36]
  wire  CAMLine_59_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_59_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_59_io_din; // @[cam.scala 81:36]
  wire  CAMLine_59_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_60_clock; // @[cam.scala 81:36]
  wire  CAMLine_60_io_we; // @[cam.scala 81:36]
  wire  CAMLine_60_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_60_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_60_io_din; // @[cam.scala 81:36]
  wire  CAMLine_60_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_61_clock; // @[cam.scala 81:36]
  wire  CAMLine_61_io_we; // @[cam.scala 81:36]
  wire  CAMLine_61_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_61_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_61_io_din; // @[cam.scala 81:36]
  wire  CAMLine_61_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_62_clock; // @[cam.scala 81:36]
  wire  CAMLine_62_io_we; // @[cam.scala 81:36]
  wire  CAMLine_62_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_62_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_62_io_din; // @[cam.scala 81:36]
  wire  CAMLine_62_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_63_clock; // @[cam.scala 81:36]
  wire  CAMLine_63_io_we; // @[cam.scala 81:36]
  wire  CAMLine_63_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_63_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_63_io_din; // @[cam.scala 81:36]
  wire  CAMLine_63_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_64_clock; // @[cam.scala 81:36]
  wire  CAMLine_64_io_we; // @[cam.scala 81:36]
  wire  CAMLine_64_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_64_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_64_io_din; // @[cam.scala 81:36]
  wire  CAMLine_64_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_65_clock; // @[cam.scala 81:36]
  wire  CAMLine_65_io_we; // @[cam.scala 81:36]
  wire  CAMLine_65_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_65_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_65_io_din; // @[cam.scala 81:36]
  wire  CAMLine_65_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_66_clock; // @[cam.scala 81:36]
  wire  CAMLine_66_io_we; // @[cam.scala 81:36]
  wire  CAMLine_66_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_66_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_66_io_din; // @[cam.scala 81:36]
  wire  CAMLine_66_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_67_clock; // @[cam.scala 81:36]
  wire  CAMLine_67_io_we; // @[cam.scala 81:36]
  wire  CAMLine_67_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_67_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_67_io_din; // @[cam.scala 81:36]
  wire  CAMLine_67_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_68_clock; // @[cam.scala 81:36]
  wire  CAMLine_68_io_we; // @[cam.scala 81:36]
  wire  CAMLine_68_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_68_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_68_io_din; // @[cam.scala 81:36]
  wire  CAMLine_68_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_69_clock; // @[cam.scala 81:36]
  wire  CAMLine_69_io_we; // @[cam.scala 81:36]
  wire  CAMLine_69_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_69_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_69_io_din; // @[cam.scala 81:36]
  wire  CAMLine_69_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_70_clock; // @[cam.scala 81:36]
  wire  CAMLine_70_io_we; // @[cam.scala 81:36]
  wire  CAMLine_70_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_70_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_70_io_din; // @[cam.scala 81:36]
  wire  CAMLine_70_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_71_clock; // @[cam.scala 81:36]
  wire  CAMLine_71_io_we; // @[cam.scala 81:36]
  wire  CAMLine_71_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_71_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_71_io_din; // @[cam.scala 81:36]
  wire  CAMLine_71_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_72_clock; // @[cam.scala 81:36]
  wire  CAMLine_72_io_we; // @[cam.scala 81:36]
  wire  CAMLine_72_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_72_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_72_io_din; // @[cam.scala 81:36]
  wire  CAMLine_72_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_73_clock; // @[cam.scala 81:36]
  wire  CAMLine_73_io_we; // @[cam.scala 81:36]
  wire  CAMLine_73_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_73_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_73_io_din; // @[cam.scala 81:36]
  wire  CAMLine_73_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_74_clock; // @[cam.scala 81:36]
  wire  CAMLine_74_io_we; // @[cam.scala 81:36]
  wire  CAMLine_74_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_74_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_74_io_din; // @[cam.scala 81:36]
  wire  CAMLine_74_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_75_clock; // @[cam.scala 81:36]
  wire  CAMLine_75_io_we; // @[cam.scala 81:36]
  wire  CAMLine_75_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_75_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_75_io_din; // @[cam.scala 81:36]
  wire  CAMLine_75_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_76_clock; // @[cam.scala 81:36]
  wire  CAMLine_76_io_we; // @[cam.scala 81:36]
  wire  CAMLine_76_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_76_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_76_io_din; // @[cam.scala 81:36]
  wire  CAMLine_76_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_77_clock; // @[cam.scala 81:36]
  wire  CAMLine_77_io_we; // @[cam.scala 81:36]
  wire  CAMLine_77_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_77_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_77_io_din; // @[cam.scala 81:36]
  wire  CAMLine_77_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_78_clock; // @[cam.scala 81:36]
  wire  CAMLine_78_io_we; // @[cam.scala 81:36]
  wire  CAMLine_78_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_78_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_78_io_din; // @[cam.scala 81:36]
  wire  CAMLine_78_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_79_clock; // @[cam.scala 81:36]
  wire  CAMLine_79_io_we; // @[cam.scala 81:36]
  wire  CAMLine_79_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_79_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_79_io_din; // @[cam.scala 81:36]
  wire  CAMLine_79_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_80_clock; // @[cam.scala 81:36]
  wire  CAMLine_80_io_we; // @[cam.scala 81:36]
  wire  CAMLine_80_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_80_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_80_io_din; // @[cam.scala 81:36]
  wire  CAMLine_80_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_81_clock; // @[cam.scala 81:36]
  wire  CAMLine_81_io_we; // @[cam.scala 81:36]
  wire  CAMLine_81_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_81_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_81_io_din; // @[cam.scala 81:36]
  wire  CAMLine_81_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_82_clock; // @[cam.scala 81:36]
  wire  CAMLine_82_io_we; // @[cam.scala 81:36]
  wire  CAMLine_82_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_82_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_82_io_din; // @[cam.scala 81:36]
  wire  CAMLine_82_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_83_clock; // @[cam.scala 81:36]
  wire  CAMLine_83_io_we; // @[cam.scala 81:36]
  wire  CAMLine_83_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_83_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_83_io_din; // @[cam.scala 81:36]
  wire  CAMLine_83_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_84_clock; // @[cam.scala 81:36]
  wire  CAMLine_84_io_we; // @[cam.scala 81:36]
  wire  CAMLine_84_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_84_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_84_io_din; // @[cam.scala 81:36]
  wire  CAMLine_84_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_85_clock; // @[cam.scala 81:36]
  wire  CAMLine_85_io_we; // @[cam.scala 81:36]
  wire  CAMLine_85_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_85_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_85_io_din; // @[cam.scala 81:36]
  wire  CAMLine_85_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_86_clock; // @[cam.scala 81:36]
  wire  CAMLine_86_io_we; // @[cam.scala 81:36]
  wire  CAMLine_86_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_86_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_86_io_din; // @[cam.scala 81:36]
  wire  CAMLine_86_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_87_clock; // @[cam.scala 81:36]
  wire  CAMLine_87_io_we; // @[cam.scala 81:36]
  wire  CAMLine_87_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_87_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_87_io_din; // @[cam.scala 81:36]
  wire  CAMLine_87_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_88_clock; // @[cam.scala 81:36]
  wire  CAMLine_88_io_we; // @[cam.scala 81:36]
  wire  CAMLine_88_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_88_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_88_io_din; // @[cam.scala 81:36]
  wire  CAMLine_88_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_89_clock; // @[cam.scala 81:36]
  wire  CAMLine_89_io_we; // @[cam.scala 81:36]
  wire  CAMLine_89_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_89_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_89_io_din; // @[cam.scala 81:36]
  wire  CAMLine_89_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_90_clock; // @[cam.scala 81:36]
  wire  CAMLine_90_io_we; // @[cam.scala 81:36]
  wire  CAMLine_90_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_90_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_90_io_din; // @[cam.scala 81:36]
  wire  CAMLine_90_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_91_clock; // @[cam.scala 81:36]
  wire  CAMLine_91_io_we; // @[cam.scala 81:36]
  wire  CAMLine_91_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_91_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_91_io_din; // @[cam.scala 81:36]
  wire  CAMLine_91_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_92_clock; // @[cam.scala 81:36]
  wire  CAMLine_92_io_we; // @[cam.scala 81:36]
  wire  CAMLine_92_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_92_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_92_io_din; // @[cam.scala 81:36]
  wire  CAMLine_92_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_93_clock; // @[cam.scala 81:36]
  wire  CAMLine_93_io_we; // @[cam.scala 81:36]
  wire  CAMLine_93_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_93_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_93_io_din; // @[cam.scala 81:36]
  wire  CAMLine_93_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_94_clock; // @[cam.scala 81:36]
  wire  CAMLine_94_io_we; // @[cam.scala 81:36]
  wire  CAMLine_94_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_94_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_94_io_din; // @[cam.scala 81:36]
  wire  CAMLine_94_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_95_clock; // @[cam.scala 81:36]
  wire  CAMLine_95_io_we; // @[cam.scala 81:36]
  wire  CAMLine_95_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_95_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_95_io_din; // @[cam.scala 81:36]
  wire  CAMLine_95_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_96_clock; // @[cam.scala 81:36]
  wire  CAMLine_96_io_we; // @[cam.scala 81:36]
  wire  CAMLine_96_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_96_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_96_io_din; // @[cam.scala 81:36]
  wire  CAMLine_96_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_97_clock; // @[cam.scala 81:36]
  wire  CAMLine_97_io_we; // @[cam.scala 81:36]
  wire  CAMLine_97_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_97_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_97_io_din; // @[cam.scala 81:36]
  wire  CAMLine_97_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_98_clock; // @[cam.scala 81:36]
  wire  CAMLine_98_io_we; // @[cam.scala 81:36]
  wire  CAMLine_98_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_98_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_98_io_din; // @[cam.scala 81:36]
  wire  CAMLine_98_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_99_clock; // @[cam.scala 81:36]
  wire  CAMLine_99_io_we; // @[cam.scala 81:36]
  wire  CAMLine_99_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_99_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_99_io_din; // @[cam.scala 81:36]
  wire  CAMLine_99_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_100_clock; // @[cam.scala 81:36]
  wire  CAMLine_100_io_we; // @[cam.scala 81:36]
  wire  CAMLine_100_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_100_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_100_io_din; // @[cam.scala 81:36]
  wire  CAMLine_100_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_101_clock; // @[cam.scala 81:36]
  wire  CAMLine_101_io_we; // @[cam.scala 81:36]
  wire  CAMLine_101_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_101_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_101_io_din; // @[cam.scala 81:36]
  wire  CAMLine_101_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_102_clock; // @[cam.scala 81:36]
  wire  CAMLine_102_io_we; // @[cam.scala 81:36]
  wire  CAMLine_102_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_102_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_102_io_din; // @[cam.scala 81:36]
  wire  CAMLine_102_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_103_clock; // @[cam.scala 81:36]
  wire  CAMLine_103_io_we; // @[cam.scala 81:36]
  wire  CAMLine_103_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_103_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_103_io_din; // @[cam.scala 81:36]
  wire  CAMLine_103_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_104_clock; // @[cam.scala 81:36]
  wire  CAMLine_104_io_we; // @[cam.scala 81:36]
  wire  CAMLine_104_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_104_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_104_io_din; // @[cam.scala 81:36]
  wire  CAMLine_104_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_105_clock; // @[cam.scala 81:36]
  wire  CAMLine_105_io_we; // @[cam.scala 81:36]
  wire  CAMLine_105_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_105_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_105_io_din; // @[cam.scala 81:36]
  wire  CAMLine_105_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_106_clock; // @[cam.scala 81:36]
  wire  CAMLine_106_io_we; // @[cam.scala 81:36]
  wire  CAMLine_106_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_106_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_106_io_din; // @[cam.scala 81:36]
  wire  CAMLine_106_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_107_clock; // @[cam.scala 81:36]
  wire  CAMLine_107_io_we; // @[cam.scala 81:36]
  wire  CAMLine_107_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_107_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_107_io_din; // @[cam.scala 81:36]
  wire  CAMLine_107_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_108_clock; // @[cam.scala 81:36]
  wire  CAMLine_108_io_we; // @[cam.scala 81:36]
  wire  CAMLine_108_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_108_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_108_io_din; // @[cam.scala 81:36]
  wire  CAMLine_108_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_109_clock; // @[cam.scala 81:36]
  wire  CAMLine_109_io_we; // @[cam.scala 81:36]
  wire  CAMLine_109_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_109_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_109_io_din; // @[cam.scala 81:36]
  wire  CAMLine_109_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_110_clock; // @[cam.scala 81:36]
  wire  CAMLine_110_io_we; // @[cam.scala 81:36]
  wire  CAMLine_110_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_110_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_110_io_din; // @[cam.scala 81:36]
  wire  CAMLine_110_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_111_clock; // @[cam.scala 81:36]
  wire  CAMLine_111_io_we; // @[cam.scala 81:36]
  wire  CAMLine_111_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_111_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_111_io_din; // @[cam.scala 81:36]
  wire  CAMLine_111_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_112_clock; // @[cam.scala 81:36]
  wire  CAMLine_112_io_we; // @[cam.scala 81:36]
  wire  CAMLine_112_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_112_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_112_io_din; // @[cam.scala 81:36]
  wire  CAMLine_112_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_113_clock; // @[cam.scala 81:36]
  wire  CAMLine_113_io_we; // @[cam.scala 81:36]
  wire  CAMLine_113_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_113_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_113_io_din; // @[cam.scala 81:36]
  wire  CAMLine_113_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_114_clock; // @[cam.scala 81:36]
  wire  CAMLine_114_io_we; // @[cam.scala 81:36]
  wire  CAMLine_114_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_114_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_114_io_din; // @[cam.scala 81:36]
  wire  CAMLine_114_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_115_clock; // @[cam.scala 81:36]
  wire  CAMLine_115_io_we; // @[cam.scala 81:36]
  wire  CAMLine_115_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_115_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_115_io_din; // @[cam.scala 81:36]
  wire  CAMLine_115_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_116_clock; // @[cam.scala 81:36]
  wire  CAMLine_116_io_we; // @[cam.scala 81:36]
  wire  CAMLine_116_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_116_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_116_io_din; // @[cam.scala 81:36]
  wire  CAMLine_116_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_117_clock; // @[cam.scala 81:36]
  wire  CAMLine_117_io_we; // @[cam.scala 81:36]
  wire  CAMLine_117_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_117_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_117_io_din; // @[cam.scala 81:36]
  wire  CAMLine_117_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_118_clock; // @[cam.scala 81:36]
  wire  CAMLine_118_io_we; // @[cam.scala 81:36]
  wire  CAMLine_118_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_118_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_118_io_din; // @[cam.scala 81:36]
  wire  CAMLine_118_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_119_clock; // @[cam.scala 81:36]
  wire  CAMLine_119_io_we; // @[cam.scala 81:36]
  wire  CAMLine_119_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_119_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_119_io_din; // @[cam.scala 81:36]
  wire  CAMLine_119_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_120_clock; // @[cam.scala 81:36]
  wire  CAMLine_120_io_we; // @[cam.scala 81:36]
  wire  CAMLine_120_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_120_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_120_io_din; // @[cam.scala 81:36]
  wire  CAMLine_120_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_121_clock; // @[cam.scala 81:36]
  wire  CAMLine_121_io_we; // @[cam.scala 81:36]
  wire  CAMLine_121_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_121_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_121_io_din; // @[cam.scala 81:36]
  wire  CAMLine_121_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_122_clock; // @[cam.scala 81:36]
  wire  CAMLine_122_io_we; // @[cam.scala 81:36]
  wire  CAMLine_122_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_122_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_122_io_din; // @[cam.scala 81:36]
  wire  CAMLine_122_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_123_clock; // @[cam.scala 81:36]
  wire  CAMLine_123_io_we; // @[cam.scala 81:36]
  wire  CAMLine_123_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_123_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_123_io_din; // @[cam.scala 81:36]
  wire  CAMLine_123_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_124_clock; // @[cam.scala 81:36]
  wire  CAMLine_124_io_we; // @[cam.scala 81:36]
  wire  CAMLine_124_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_124_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_124_io_din; // @[cam.scala 81:36]
  wire  CAMLine_124_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_125_clock; // @[cam.scala 81:36]
  wire  CAMLine_125_io_we; // @[cam.scala 81:36]
  wire  CAMLine_125_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_125_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_125_io_din; // @[cam.scala 81:36]
  wire  CAMLine_125_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_126_clock; // @[cam.scala 81:36]
  wire  CAMLine_126_io_we; // @[cam.scala 81:36]
  wire  CAMLine_126_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_126_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_126_io_din; // @[cam.scala 81:36]
  wire  CAMLine_126_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_127_clock; // @[cam.scala 81:36]
  wire  CAMLine_127_io_we; // @[cam.scala 81:36]
  wire  CAMLine_127_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_127_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_127_io_din; // @[cam.scala 81:36]
  wire  CAMLine_127_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_128_clock; // @[cam.scala 81:36]
  wire  CAMLine_128_io_we; // @[cam.scala 81:36]
  wire  CAMLine_128_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_128_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_128_io_din; // @[cam.scala 81:36]
  wire  CAMLine_128_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_129_clock; // @[cam.scala 81:36]
  wire  CAMLine_129_io_we; // @[cam.scala 81:36]
  wire  CAMLine_129_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_129_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_129_io_din; // @[cam.scala 81:36]
  wire  CAMLine_129_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_130_clock; // @[cam.scala 81:36]
  wire  CAMLine_130_io_we; // @[cam.scala 81:36]
  wire  CAMLine_130_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_130_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_130_io_din; // @[cam.scala 81:36]
  wire  CAMLine_130_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_131_clock; // @[cam.scala 81:36]
  wire  CAMLine_131_io_we; // @[cam.scala 81:36]
  wire  CAMLine_131_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_131_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_131_io_din; // @[cam.scala 81:36]
  wire  CAMLine_131_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_132_clock; // @[cam.scala 81:36]
  wire  CAMLine_132_io_we; // @[cam.scala 81:36]
  wire  CAMLine_132_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_132_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_132_io_din; // @[cam.scala 81:36]
  wire  CAMLine_132_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_133_clock; // @[cam.scala 81:36]
  wire  CAMLine_133_io_we; // @[cam.scala 81:36]
  wire  CAMLine_133_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_133_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_133_io_din; // @[cam.scala 81:36]
  wire  CAMLine_133_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_134_clock; // @[cam.scala 81:36]
  wire  CAMLine_134_io_we; // @[cam.scala 81:36]
  wire  CAMLine_134_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_134_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_134_io_din; // @[cam.scala 81:36]
  wire  CAMLine_134_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_135_clock; // @[cam.scala 81:36]
  wire  CAMLine_135_io_we; // @[cam.scala 81:36]
  wire  CAMLine_135_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_135_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_135_io_din; // @[cam.scala 81:36]
  wire  CAMLine_135_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_136_clock; // @[cam.scala 81:36]
  wire  CAMLine_136_io_we; // @[cam.scala 81:36]
  wire  CAMLine_136_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_136_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_136_io_din; // @[cam.scala 81:36]
  wire  CAMLine_136_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_137_clock; // @[cam.scala 81:36]
  wire  CAMLine_137_io_we; // @[cam.scala 81:36]
  wire  CAMLine_137_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_137_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_137_io_din; // @[cam.scala 81:36]
  wire  CAMLine_137_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_138_clock; // @[cam.scala 81:36]
  wire  CAMLine_138_io_we; // @[cam.scala 81:36]
  wire  CAMLine_138_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_138_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_138_io_din; // @[cam.scala 81:36]
  wire  CAMLine_138_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_139_clock; // @[cam.scala 81:36]
  wire  CAMLine_139_io_we; // @[cam.scala 81:36]
  wire  CAMLine_139_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_139_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_139_io_din; // @[cam.scala 81:36]
  wire  CAMLine_139_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_140_clock; // @[cam.scala 81:36]
  wire  CAMLine_140_io_we; // @[cam.scala 81:36]
  wire  CAMLine_140_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_140_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_140_io_din; // @[cam.scala 81:36]
  wire  CAMLine_140_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_141_clock; // @[cam.scala 81:36]
  wire  CAMLine_141_io_we; // @[cam.scala 81:36]
  wire  CAMLine_141_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_141_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_141_io_din; // @[cam.scala 81:36]
  wire  CAMLine_141_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_142_clock; // @[cam.scala 81:36]
  wire  CAMLine_142_io_we; // @[cam.scala 81:36]
  wire  CAMLine_142_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_142_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_142_io_din; // @[cam.scala 81:36]
  wire  CAMLine_142_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_143_clock; // @[cam.scala 81:36]
  wire  CAMLine_143_io_we; // @[cam.scala 81:36]
  wire  CAMLine_143_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_143_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_143_io_din; // @[cam.scala 81:36]
  wire  CAMLine_143_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_144_clock; // @[cam.scala 81:36]
  wire  CAMLine_144_io_we; // @[cam.scala 81:36]
  wire  CAMLine_144_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_144_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_144_io_din; // @[cam.scala 81:36]
  wire  CAMLine_144_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_145_clock; // @[cam.scala 81:36]
  wire  CAMLine_145_io_we; // @[cam.scala 81:36]
  wire  CAMLine_145_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_145_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_145_io_din; // @[cam.scala 81:36]
  wire  CAMLine_145_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_146_clock; // @[cam.scala 81:36]
  wire  CAMLine_146_io_we; // @[cam.scala 81:36]
  wire  CAMLine_146_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_146_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_146_io_din; // @[cam.scala 81:36]
  wire  CAMLine_146_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_147_clock; // @[cam.scala 81:36]
  wire  CAMLine_147_io_we; // @[cam.scala 81:36]
  wire  CAMLine_147_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_147_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_147_io_din; // @[cam.scala 81:36]
  wire  CAMLine_147_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_148_clock; // @[cam.scala 81:36]
  wire  CAMLine_148_io_we; // @[cam.scala 81:36]
  wire  CAMLine_148_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_148_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_148_io_din; // @[cam.scala 81:36]
  wire  CAMLine_148_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_149_clock; // @[cam.scala 81:36]
  wire  CAMLine_149_io_we; // @[cam.scala 81:36]
  wire  CAMLine_149_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_149_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_149_io_din; // @[cam.scala 81:36]
  wire  CAMLine_149_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_150_clock; // @[cam.scala 81:36]
  wire  CAMLine_150_io_we; // @[cam.scala 81:36]
  wire  CAMLine_150_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_150_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_150_io_din; // @[cam.scala 81:36]
  wire  CAMLine_150_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_151_clock; // @[cam.scala 81:36]
  wire  CAMLine_151_io_we; // @[cam.scala 81:36]
  wire  CAMLine_151_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_151_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_151_io_din; // @[cam.scala 81:36]
  wire  CAMLine_151_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_152_clock; // @[cam.scala 81:36]
  wire  CAMLine_152_io_we; // @[cam.scala 81:36]
  wire  CAMLine_152_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_152_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_152_io_din; // @[cam.scala 81:36]
  wire  CAMLine_152_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_153_clock; // @[cam.scala 81:36]
  wire  CAMLine_153_io_we; // @[cam.scala 81:36]
  wire  CAMLine_153_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_153_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_153_io_din; // @[cam.scala 81:36]
  wire  CAMLine_153_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_154_clock; // @[cam.scala 81:36]
  wire  CAMLine_154_io_we; // @[cam.scala 81:36]
  wire  CAMLine_154_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_154_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_154_io_din; // @[cam.scala 81:36]
  wire  CAMLine_154_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_155_clock; // @[cam.scala 81:36]
  wire  CAMLine_155_io_we; // @[cam.scala 81:36]
  wire  CAMLine_155_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_155_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_155_io_din; // @[cam.scala 81:36]
  wire  CAMLine_155_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_156_clock; // @[cam.scala 81:36]
  wire  CAMLine_156_io_we; // @[cam.scala 81:36]
  wire  CAMLine_156_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_156_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_156_io_din; // @[cam.scala 81:36]
  wire  CAMLine_156_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_157_clock; // @[cam.scala 81:36]
  wire  CAMLine_157_io_we; // @[cam.scala 81:36]
  wire  CAMLine_157_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_157_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_157_io_din; // @[cam.scala 81:36]
  wire  CAMLine_157_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_158_clock; // @[cam.scala 81:36]
  wire  CAMLine_158_io_we; // @[cam.scala 81:36]
  wire  CAMLine_158_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_158_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_158_io_din; // @[cam.scala 81:36]
  wire  CAMLine_158_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_159_clock; // @[cam.scala 81:36]
  wire  CAMLine_159_io_we; // @[cam.scala 81:36]
  wire  CAMLine_159_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_159_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_159_io_din; // @[cam.scala 81:36]
  wire  CAMLine_159_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_160_clock; // @[cam.scala 81:36]
  wire  CAMLine_160_io_we; // @[cam.scala 81:36]
  wire  CAMLine_160_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_160_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_160_io_din; // @[cam.scala 81:36]
  wire  CAMLine_160_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_161_clock; // @[cam.scala 81:36]
  wire  CAMLine_161_io_we; // @[cam.scala 81:36]
  wire  CAMLine_161_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_161_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_161_io_din; // @[cam.scala 81:36]
  wire  CAMLine_161_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_162_clock; // @[cam.scala 81:36]
  wire  CAMLine_162_io_we; // @[cam.scala 81:36]
  wire  CAMLine_162_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_162_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_162_io_din; // @[cam.scala 81:36]
  wire  CAMLine_162_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_163_clock; // @[cam.scala 81:36]
  wire  CAMLine_163_io_we; // @[cam.scala 81:36]
  wire  CAMLine_163_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_163_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_163_io_din; // @[cam.scala 81:36]
  wire  CAMLine_163_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_164_clock; // @[cam.scala 81:36]
  wire  CAMLine_164_io_we; // @[cam.scala 81:36]
  wire  CAMLine_164_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_164_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_164_io_din; // @[cam.scala 81:36]
  wire  CAMLine_164_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_165_clock; // @[cam.scala 81:36]
  wire  CAMLine_165_io_we; // @[cam.scala 81:36]
  wire  CAMLine_165_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_165_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_165_io_din; // @[cam.scala 81:36]
  wire  CAMLine_165_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_166_clock; // @[cam.scala 81:36]
  wire  CAMLine_166_io_we; // @[cam.scala 81:36]
  wire  CAMLine_166_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_166_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_166_io_din; // @[cam.scala 81:36]
  wire  CAMLine_166_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_167_clock; // @[cam.scala 81:36]
  wire  CAMLine_167_io_we; // @[cam.scala 81:36]
  wire  CAMLine_167_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_167_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_167_io_din; // @[cam.scala 81:36]
  wire  CAMLine_167_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_168_clock; // @[cam.scala 81:36]
  wire  CAMLine_168_io_we; // @[cam.scala 81:36]
  wire  CAMLine_168_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_168_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_168_io_din; // @[cam.scala 81:36]
  wire  CAMLine_168_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_169_clock; // @[cam.scala 81:36]
  wire  CAMLine_169_io_we; // @[cam.scala 81:36]
  wire  CAMLine_169_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_169_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_169_io_din; // @[cam.scala 81:36]
  wire  CAMLine_169_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_170_clock; // @[cam.scala 81:36]
  wire  CAMLine_170_io_we; // @[cam.scala 81:36]
  wire  CAMLine_170_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_170_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_170_io_din; // @[cam.scala 81:36]
  wire  CAMLine_170_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_171_clock; // @[cam.scala 81:36]
  wire  CAMLine_171_io_we; // @[cam.scala 81:36]
  wire  CAMLine_171_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_171_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_171_io_din; // @[cam.scala 81:36]
  wire  CAMLine_171_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_172_clock; // @[cam.scala 81:36]
  wire  CAMLine_172_io_we; // @[cam.scala 81:36]
  wire  CAMLine_172_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_172_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_172_io_din; // @[cam.scala 81:36]
  wire  CAMLine_172_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_173_clock; // @[cam.scala 81:36]
  wire  CAMLine_173_io_we; // @[cam.scala 81:36]
  wire  CAMLine_173_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_173_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_173_io_din; // @[cam.scala 81:36]
  wire  CAMLine_173_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_174_clock; // @[cam.scala 81:36]
  wire  CAMLine_174_io_we; // @[cam.scala 81:36]
  wire  CAMLine_174_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_174_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_174_io_din; // @[cam.scala 81:36]
  wire  CAMLine_174_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_175_clock; // @[cam.scala 81:36]
  wire  CAMLine_175_io_we; // @[cam.scala 81:36]
  wire  CAMLine_175_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_175_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_175_io_din; // @[cam.scala 81:36]
  wire  CAMLine_175_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_176_clock; // @[cam.scala 81:36]
  wire  CAMLine_176_io_we; // @[cam.scala 81:36]
  wire  CAMLine_176_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_176_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_176_io_din; // @[cam.scala 81:36]
  wire  CAMLine_176_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_177_clock; // @[cam.scala 81:36]
  wire  CAMLine_177_io_we; // @[cam.scala 81:36]
  wire  CAMLine_177_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_177_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_177_io_din; // @[cam.scala 81:36]
  wire  CAMLine_177_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_178_clock; // @[cam.scala 81:36]
  wire  CAMLine_178_io_we; // @[cam.scala 81:36]
  wire  CAMLine_178_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_178_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_178_io_din; // @[cam.scala 81:36]
  wire  CAMLine_178_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_179_clock; // @[cam.scala 81:36]
  wire  CAMLine_179_io_we; // @[cam.scala 81:36]
  wire  CAMLine_179_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_179_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_179_io_din; // @[cam.scala 81:36]
  wire  CAMLine_179_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_180_clock; // @[cam.scala 81:36]
  wire  CAMLine_180_io_we; // @[cam.scala 81:36]
  wire  CAMLine_180_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_180_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_180_io_din; // @[cam.scala 81:36]
  wire  CAMLine_180_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_181_clock; // @[cam.scala 81:36]
  wire  CAMLine_181_io_we; // @[cam.scala 81:36]
  wire  CAMLine_181_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_181_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_181_io_din; // @[cam.scala 81:36]
  wire  CAMLine_181_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_182_clock; // @[cam.scala 81:36]
  wire  CAMLine_182_io_we; // @[cam.scala 81:36]
  wire  CAMLine_182_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_182_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_182_io_din; // @[cam.scala 81:36]
  wire  CAMLine_182_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_183_clock; // @[cam.scala 81:36]
  wire  CAMLine_183_io_we; // @[cam.scala 81:36]
  wire  CAMLine_183_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_183_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_183_io_din; // @[cam.scala 81:36]
  wire  CAMLine_183_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_184_clock; // @[cam.scala 81:36]
  wire  CAMLine_184_io_we; // @[cam.scala 81:36]
  wire  CAMLine_184_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_184_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_184_io_din; // @[cam.scala 81:36]
  wire  CAMLine_184_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_185_clock; // @[cam.scala 81:36]
  wire  CAMLine_185_io_we; // @[cam.scala 81:36]
  wire  CAMLine_185_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_185_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_185_io_din; // @[cam.scala 81:36]
  wire  CAMLine_185_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_186_clock; // @[cam.scala 81:36]
  wire  CAMLine_186_io_we; // @[cam.scala 81:36]
  wire  CAMLine_186_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_186_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_186_io_din; // @[cam.scala 81:36]
  wire  CAMLine_186_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_187_clock; // @[cam.scala 81:36]
  wire  CAMLine_187_io_we; // @[cam.scala 81:36]
  wire  CAMLine_187_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_187_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_187_io_din; // @[cam.scala 81:36]
  wire  CAMLine_187_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_188_clock; // @[cam.scala 81:36]
  wire  CAMLine_188_io_we; // @[cam.scala 81:36]
  wire  CAMLine_188_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_188_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_188_io_din; // @[cam.scala 81:36]
  wire  CAMLine_188_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_189_clock; // @[cam.scala 81:36]
  wire  CAMLine_189_io_we; // @[cam.scala 81:36]
  wire  CAMLine_189_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_189_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_189_io_din; // @[cam.scala 81:36]
  wire  CAMLine_189_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_190_clock; // @[cam.scala 81:36]
  wire  CAMLine_190_io_we; // @[cam.scala 81:36]
  wire  CAMLine_190_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_190_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_190_io_din; // @[cam.scala 81:36]
  wire  CAMLine_190_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_191_clock; // @[cam.scala 81:36]
  wire  CAMLine_191_io_we; // @[cam.scala 81:36]
  wire  CAMLine_191_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_191_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_191_io_din; // @[cam.scala 81:36]
  wire  CAMLine_191_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_192_clock; // @[cam.scala 81:36]
  wire  CAMLine_192_io_we; // @[cam.scala 81:36]
  wire  CAMLine_192_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_192_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_192_io_din; // @[cam.scala 81:36]
  wire  CAMLine_192_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_193_clock; // @[cam.scala 81:36]
  wire  CAMLine_193_io_we; // @[cam.scala 81:36]
  wire  CAMLine_193_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_193_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_193_io_din; // @[cam.scala 81:36]
  wire  CAMLine_193_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_194_clock; // @[cam.scala 81:36]
  wire  CAMLine_194_io_we; // @[cam.scala 81:36]
  wire  CAMLine_194_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_194_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_194_io_din; // @[cam.scala 81:36]
  wire  CAMLine_194_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_195_clock; // @[cam.scala 81:36]
  wire  CAMLine_195_io_we; // @[cam.scala 81:36]
  wire  CAMLine_195_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_195_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_195_io_din; // @[cam.scala 81:36]
  wire  CAMLine_195_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_196_clock; // @[cam.scala 81:36]
  wire  CAMLine_196_io_we; // @[cam.scala 81:36]
  wire  CAMLine_196_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_196_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_196_io_din; // @[cam.scala 81:36]
  wire  CAMLine_196_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_197_clock; // @[cam.scala 81:36]
  wire  CAMLine_197_io_we; // @[cam.scala 81:36]
  wire  CAMLine_197_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_197_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_197_io_din; // @[cam.scala 81:36]
  wire  CAMLine_197_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_198_clock; // @[cam.scala 81:36]
  wire  CAMLine_198_io_we; // @[cam.scala 81:36]
  wire  CAMLine_198_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_198_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_198_io_din; // @[cam.scala 81:36]
  wire  CAMLine_198_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_199_clock; // @[cam.scala 81:36]
  wire  CAMLine_199_io_we; // @[cam.scala 81:36]
  wire  CAMLine_199_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_199_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_199_io_din; // @[cam.scala 81:36]
  wire  CAMLine_199_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_200_clock; // @[cam.scala 81:36]
  wire  CAMLine_200_io_we; // @[cam.scala 81:36]
  wire  CAMLine_200_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_200_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_200_io_din; // @[cam.scala 81:36]
  wire  CAMLine_200_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_201_clock; // @[cam.scala 81:36]
  wire  CAMLine_201_io_we; // @[cam.scala 81:36]
  wire  CAMLine_201_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_201_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_201_io_din; // @[cam.scala 81:36]
  wire  CAMLine_201_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_202_clock; // @[cam.scala 81:36]
  wire  CAMLine_202_io_we; // @[cam.scala 81:36]
  wire  CAMLine_202_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_202_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_202_io_din; // @[cam.scala 81:36]
  wire  CAMLine_202_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_203_clock; // @[cam.scala 81:36]
  wire  CAMLine_203_io_we; // @[cam.scala 81:36]
  wire  CAMLine_203_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_203_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_203_io_din; // @[cam.scala 81:36]
  wire  CAMLine_203_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_204_clock; // @[cam.scala 81:36]
  wire  CAMLine_204_io_we; // @[cam.scala 81:36]
  wire  CAMLine_204_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_204_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_204_io_din; // @[cam.scala 81:36]
  wire  CAMLine_204_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_205_clock; // @[cam.scala 81:36]
  wire  CAMLine_205_io_we; // @[cam.scala 81:36]
  wire  CAMLine_205_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_205_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_205_io_din; // @[cam.scala 81:36]
  wire  CAMLine_205_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_206_clock; // @[cam.scala 81:36]
  wire  CAMLine_206_io_we; // @[cam.scala 81:36]
  wire  CAMLine_206_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_206_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_206_io_din; // @[cam.scala 81:36]
  wire  CAMLine_206_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_207_clock; // @[cam.scala 81:36]
  wire  CAMLine_207_io_we; // @[cam.scala 81:36]
  wire  CAMLine_207_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_207_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_207_io_din; // @[cam.scala 81:36]
  wire  CAMLine_207_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_208_clock; // @[cam.scala 81:36]
  wire  CAMLine_208_io_we; // @[cam.scala 81:36]
  wire  CAMLine_208_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_208_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_208_io_din; // @[cam.scala 81:36]
  wire  CAMLine_208_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_209_clock; // @[cam.scala 81:36]
  wire  CAMLine_209_io_we; // @[cam.scala 81:36]
  wire  CAMLine_209_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_209_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_209_io_din; // @[cam.scala 81:36]
  wire  CAMLine_209_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_210_clock; // @[cam.scala 81:36]
  wire  CAMLine_210_io_we; // @[cam.scala 81:36]
  wire  CAMLine_210_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_210_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_210_io_din; // @[cam.scala 81:36]
  wire  CAMLine_210_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_211_clock; // @[cam.scala 81:36]
  wire  CAMLine_211_io_we; // @[cam.scala 81:36]
  wire  CAMLine_211_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_211_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_211_io_din; // @[cam.scala 81:36]
  wire  CAMLine_211_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_212_clock; // @[cam.scala 81:36]
  wire  CAMLine_212_io_we; // @[cam.scala 81:36]
  wire  CAMLine_212_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_212_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_212_io_din; // @[cam.scala 81:36]
  wire  CAMLine_212_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_213_clock; // @[cam.scala 81:36]
  wire  CAMLine_213_io_we; // @[cam.scala 81:36]
  wire  CAMLine_213_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_213_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_213_io_din; // @[cam.scala 81:36]
  wire  CAMLine_213_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_214_clock; // @[cam.scala 81:36]
  wire  CAMLine_214_io_we; // @[cam.scala 81:36]
  wire  CAMLine_214_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_214_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_214_io_din; // @[cam.scala 81:36]
  wire  CAMLine_214_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_215_clock; // @[cam.scala 81:36]
  wire  CAMLine_215_io_we; // @[cam.scala 81:36]
  wire  CAMLine_215_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_215_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_215_io_din; // @[cam.scala 81:36]
  wire  CAMLine_215_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_216_clock; // @[cam.scala 81:36]
  wire  CAMLine_216_io_we; // @[cam.scala 81:36]
  wire  CAMLine_216_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_216_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_216_io_din; // @[cam.scala 81:36]
  wire  CAMLine_216_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_217_clock; // @[cam.scala 81:36]
  wire  CAMLine_217_io_we; // @[cam.scala 81:36]
  wire  CAMLine_217_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_217_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_217_io_din; // @[cam.scala 81:36]
  wire  CAMLine_217_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_218_clock; // @[cam.scala 81:36]
  wire  CAMLine_218_io_we; // @[cam.scala 81:36]
  wire  CAMLine_218_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_218_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_218_io_din; // @[cam.scala 81:36]
  wire  CAMLine_218_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_219_clock; // @[cam.scala 81:36]
  wire  CAMLine_219_io_we; // @[cam.scala 81:36]
  wire  CAMLine_219_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_219_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_219_io_din; // @[cam.scala 81:36]
  wire  CAMLine_219_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_220_clock; // @[cam.scala 81:36]
  wire  CAMLine_220_io_we; // @[cam.scala 81:36]
  wire  CAMLine_220_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_220_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_220_io_din; // @[cam.scala 81:36]
  wire  CAMLine_220_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_221_clock; // @[cam.scala 81:36]
  wire  CAMLine_221_io_we; // @[cam.scala 81:36]
  wire  CAMLine_221_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_221_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_221_io_din; // @[cam.scala 81:36]
  wire  CAMLine_221_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_222_clock; // @[cam.scala 81:36]
  wire  CAMLine_222_io_we; // @[cam.scala 81:36]
  wire  CAMLine_222_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_222_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_222_io_din; // @[cam.scala 81:36]
  wire  CAMLine_222_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_223_clock; // @[cam.scala 81:36]
  wire  CAMLine_223_io_we; // @[cam.scala 81:36]
  wire  CAMLine_223_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_223_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_223_io_din; // @[cam.scala 81:36]
  wire  CAMLine_223_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_224_clock; // @[cam.scala 81:36]
  wire  CAMLine_224_io_we; // @[cam.scala 81:36]
  wire  CAMLine_224_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_224_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_224_io_din; // @[cam.scala 81:36]
  wire  CAMLine_224_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_225_clock; // @[cam.scala 81:36]
  wire  CAMLine_225_io_we; // @[cam.scala 81:36]
  wire  CAMLine_225_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_225_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_225_io_din; // @[cam.scala 81:36]
  wire  CAMLine_225_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_226_clock; // @[cam.scala 81:36]
  wire  CAMLine_226_io_we; // @[cam.scala 81:36]
  wire  CAMLine_226_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_226_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_226_io_din; // @[cam.scala 81:36]
  wire  CAMLine_226_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_227_clock; // @[cam.scala 81:36]
  wire  CAMLine_227_io_we; // @[cam.scala 81:36]
  wire  CAMLine_227_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_227_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_227_io_din; // @[cam.scala 81:36]
  wire  CAMLine_227_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_228_clock; // @[cam.scala 81:36]
  wire  CAMLine_228_io_we; // @[cam.scala 81:36]
  wire  CAMLine_228_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_228_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_228_io_din; // @[cam.scala 81:36]
  wire  CAMLine_228_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_229_clock; // @[cam.scala 81:36]
  wire  CAMLine_229_io_we; // @[cam.scala 81:36]
  wire  CAMLine_229_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_229_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_229_io_din; // @[cam.scala 81:36]
  wire  CAMLine_229_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_230_clock; // @[cam.scala 81:36]
  wire  CAMLine_230_io_we; // @[cam.scala 81:36]
  wire  CAMLine_230_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_230_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_230_io_din; // @[cam.scala 81:36]
  wire  CAMLine_230_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_231_clock; // @[cam.scala 81:36]
  wire  CAMLine_231_io_we; // @[cam.scala 81:36]
  wire  CAMLine_231_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_231_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_231_io_din; // @[cam.scala 81:36]
  wire  CAMLine_231_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_232_clock; // @[cam.scala 81:36]
  wire  CAMLine_232_io_we; // @[cam.scala 81:36]
  wire  CAMLine_232_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_232_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_232_io_din; // @[cam.scala 81:36]
  wire  CAMLine_232_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_233_clock; // @[cam.scala 81:36]
  wire  CAMLine_233_io_we; // @[cam.scala 81:36]
  wire  CAMLine_233_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_233_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_233_io_din; // @[cam.scala 81:36]
  wire  CAMLine_233_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_234_clock; // @[cam.scala 81:36]
  wire  CAMLine_234_io_we; // @[cam.scala 81:36]
  wire  CAMLine_234_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_234_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_234_io_din; // @[cam.scala 81:36]
  wire  CAMLine_234_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_235_clock; // @[cam.scala 81:36]
  wire  CAMLine_235_io_we; // @[cam.scala 81:36]
  wire  CAMLine_235_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_235_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_235_io_din; // @[cam.scala 81:36]
  wire  CAMLine_235_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_236_clock; // @[cam.scala 81:36]
  wire  CAMLine_236_io_we; // @[cam.scala 81:36]
  wire  CAMLine_236_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_236_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_236_io_din; // @[cam.scala 81:36]
  wire  CAMLine_236_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_237_clock; // @[cam.scala 81:36]
  wire  CAMLine_237_io_we; // @[cam.scala 81:36]
  wire  CAMLine_237_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_237_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_237_io_din; // @[cam.scala 81:36]
  wire  CAMLine_237_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_238_clock; // @[cam.scala 81:36]
  wire  CAMLine_238_io_we; // @[cam.scala 81:36]
  wire  CAMLine_238_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_238_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_238_io_din; // @[cam.scala 81:36]
  wire  CAMLine_238_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_239_clock; // @[cam.scala 81:36]
  wire  CAMLine_239_io_we; // @[cam.scala 81:36]
  wire  CAMLine_239_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_239_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_239_io_din; // @[cam.scala 81:36]
  wire  CAMLine_239_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_240_clock; // @[cam.scala 81:36]
  wire  CAMLine_240_io_we; // @[cam.scala 81:36]
  wire  CAMLine_240_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_240_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_240_io_din; // @[cam.scala 81:36]
  wire  CAMLine_240_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_241_clock; // @[cam.scala 81:36]
  wire  CAMLine_241_io_we; // @[cam.scala 81:36]
  wire  CAMLine_241_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_241_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_241_io_din; // @[cam.scala 81:36]
  wire  CAMLine_241_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_242_clock; // @[cam.scala 81:36]
  wire  CAMLine_242_io_we; // @[cam.scala 81:36]
  wire  CAMLine_242_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_242_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_242_io_din; // @[cam.scala 81:36]
  wire  CAMLine_242_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_243_clock; // @[cam.scala 81:36]
  wire  CAMLine_243_io_we; // @[cam.scala 81:36]
  wire  CAMLine_243_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_243_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_243_io_din; // @[cam.scala 81:36]
  wire  CAMLine_243_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_244_clock; // @[cam.scala 81:36]
  wire  CAMLine_244_io_we; // @[cam.scala 81:36]
  wire  CAMLine_244_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_244_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_244_io_din; // @[cam.scala 81:36]
  wire  CAMLine_244_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_245_clock; // @[cam.scala 81:36]
  wire  CAMLine_245_io_we; // @[cam.scala 81:36]
  wire  CAMLine_245_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_245_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_245_io_din; // @[cam.scala 81:36]
  wire  CAMLine_245_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_246_clock; // @[cam.scala 81:36]
  wire  CAMLine_246_io_we; // @[cam.scala 81:36]
  wire  CAMLine_246_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_246_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_246_io_din; // @[cam.scala 81:36]
  wire  CAMLine_246_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_247_clock; // @[cam.scala 81:36]
  wire  CAMLine_247_io_we; // @[cam.scala 81:36]
  wire  CAMLine_247_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_247_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_247_io_din; // @[cam.scala 81:36]
  wire  CAMLine_247_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_248_clock; // @[cam.scala 81:36]
  wire  CAMLine_248_io_we; // @[cam.scala 81:36]
  wire  CAMLine_248_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_248_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_248_io_din; // @[cam.scala 81:36]
  wire  CAMLine_248_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_249_clock; // @[cam.scala 81:36]
  wire  CAMLine_249_io_we; // @[cam.scala 81:36]
  wire  CAMLine_249_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_249_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_249_io_din; // @[cam.scala 81:36]
  wire  CAMLine_249_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_250_clock; // @[cam.scala 81:36]
  wire  CAMLine_250_io_we; // @[cam.scala 81:36]
  wire  CAMLine_250_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_250_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_250_io_din; // @[cam.scala 81:36]
  wire  CAMLine_250_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_251_clock; // @[cam.scala 81:36]
  wire  CAMLine_251_io_we; // @[cam.scala 81:36]
  wire  CAMLine_251_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_251_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_251_io_din; // @[cam.scala 81:36]
  wire  CAMLine_251_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_252_clock; // @[cam.scala 81:36]
  wire  CAMLine_252_io_we; // @[cam.scala 81:36]
  wire  CAMLine_252_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_252_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_252_io_din; // @[cam.scala 81:36]
  wire  CAMLine_252_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_253_clock; // @[cam.scala 81:36]
  wire  CAMLine_253_io_we; // @[cam.scala 81:36]
  wire  CAMLine_253_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_253_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_253_io_din; // @[cam.scala 81:36]
  wire  CAMLine_253_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_254_clock; // @[cam.scala 81:36]
  wire  CAMLine_254_io_we; // @[cam.scala 81:36]
  wire  CAMLine_254_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_254_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_254_io_din; // @[cam.scala 81:36]
  wire  CAMLine_254_io_hit; // @[cam.scala 81:36]
  wire  CAMLine_255_clock; // @[cam.scala 81:36]
  wire  CAMLine_255_io_we; // @[cam.scala 81:36]
  wire  CAMLine_255_io_wi; // @[cam.scala 81:36]
  wire [255:0] CAMLine_255_io_key; // @[cam.scala 81:36]
  wire [255:0] CAMLine_255_io_din; // @[cam.scala 81:36]
  wire  CAMLine_255_io_hit; // @[cam.scala 81:36]
  wire  _io_hit_T_29 = CAMLine_io_hit | CAMLine_1_io_hit | CAMLine_2_io_hit | CAMLine_3_io_hit | CAMLine_4_io_hit |
    CAMLine_5_io_hit | CAMLine_6_io_hit | CAMLine_7_io_hit | CAMLine_8_io_hit | CAMLine_9_io_hit | CAMLine_10_io_hit |
    CAMLine_11_io_hit | CAMLine_12_io_hit | CAMLine_13_io_hit | CAMLine_14_io_hit | CAMLine_15_io_hit |
    CAMLine_16_io_hit | CAMLine_17_io_hit | CAMLine_18_io_hit | CAMLine_19_io_hit | CAMLine_20_io_hit |
    CAMLine_21_io_hit | CAMLine_22_io_hit | CAMLine_23_io_hit | CAMLine_24_io_hit | CAMLine_25_io_hit |
    CAMLine_26_io_hit | CAMLine_27_io_hit | CAMLine_28_io_hit | CAMLine_29_io_hit | CAMLine_30_io_hit; // @[cam.scala 93:27]
  wire  _io_hit_T_59 = _io_hit_T_29 | CAMLine_31_io_hit | CAMLine_32_io_hit | CAMLine_33_io_hit | CAMLine_34_io_hit |
    CAMLine_35_io_hit | CAMLine_36_io_hit | CAMLine_37_io_hit | CAMLine_38_io_hit | CAMLine_39_io_hit |
    CAMLine_40_io_hit | CAMLine_41_io_hit | CAMLine_42_io_hit | CAMLine_43_io_hit | CAMLine_44_io_hit |
    CAMLine_45_io_hit | CAMLine_46_io_hit | CAMLine_47_io_hit | CAMLine_48_io_hit | CAMLine_49_io_hit |
    CAMLine_50_io_hit | CAMLine_51_io_hit | CAMLine_52_io_hit | CAMLine_53_io_hit | CAMLine_54_io_hit |
    CAMLine_55_io_hit | CAMLine_56_io_hit | CAMLine_57_io_hit | CAMLine_58_io_hit | CAMLine_59_io_hit |
    CAMLine_60_io_hit; // @[cam.scala 93:27]
  wire  _io_hit_T_89 = _io_hit_T_59 | CAMLine_61_io_hit | CAMLine_62_io_hit | CAMLine_63_io_hit | CAMLine_64_io_hit |
    CAMLine_65_io_hit | CAMLine_66_io_hit | CAMLine_67_io_hit | CAMLine_68_io_hit | CAMLine_69_io_hit |
    CAMLine_70_io_hit | CAMLine_71_io_hit | CAMLine_72_io_hit | CAMLine_73_io_hit | CAMLine_74_io_hit |
    CAMLine_75_io_hit | CAMLine_76_io_hit | CAMLine_77_io_hit | CAMLine_78_io_hit | CAMLine_79_io_hit |
    CAMLine_80_io_hit | CAMLine_81_io_hit | CAMLine_82_io_hit | CAMLine_83_io_hit | CAMLine_84_io_hit |
    CAMLine_85_io_hit | CAMLine_86_io_hit | CAMLine_87_io_hit | CAMLine_88_io_hit | CAMLine_89_io_hit |
    CAMLine_90_io_hit; // @[cam.scala 93:27]
  wire  _io_hit_T_119 = _io_hit_T_89 | CAMLine_91_io_hit | CAMLine_92_io_hit | CAMLine_93_io_hit | CAMLine_94_io_hit |
    CAMLine_95_io_hit | CAMLine_96_io_hit | CAMLine_97_io_hit | CAMLine_98_io_hit | CAMLine_99_io_hit |
    CAMLine_100_io_hit | CAMLine_101_io_hit | CAMLine_102_io_hit | CAMLine_103_io_hit | CAMLine_104_io_hit |
    CAMLine_105_io_hit | CAMLine_106_io_hit | CAMLine_107_io_hit | CAMLine_108_io_hit | CAMLine_109_io_hit |
    CAMLine_110_io_hit | CAMLine_111_io_hit | CAMLine_112_io_hit | CAMLine_113_io_hit | CAMLine_114_io_hit |
    CAMLine_115_io_hit | CAMLine_116_io_hit | CAMLine_117_io_hit | CAMLine_118_io_hit | CAMLine_119_io_hit |
    CAMLine_120_io_hit; // @[cam.scala 93:27]
  wire  _io_hit_T_149 = _io_hit_T_119 | CAMLine_121_io_hit | CAMLine_122_io_hit | CAMLine_123_io_hit |
    CAMLine_124_io_hit | CAMLine_125_io_hit | CAMLine_126_io_hit | CAMLine_127_io_hit | CAMLine_128_io_hit |
    CAMLine_129_io_hit | CAMLine_130_io_hit | CAMLine_131_io_hit | CAMLine_132_io_hit | CAMLine_133_io_hit |
    CAMLine_134_io_hit | CAMLine_135_io_hit | CAMLine_136_io_hit | CAMLine_137_io_hit | CAMLine_138_io_hit |
    CAMLine_139_io_hit | CAMLine_140_io_hit | CAMLine_141_io_hit | CAMLine_142_io_hit | CAMLine_143_io_hit |
    CAMLine_144_io_hit | CAMLine_145_io_hit | CAMLine_146_io_hit | CAMLine_147_io_hit | CAMLine_148_io_hit |
    CAMLine_149_io_hit | CAMLine_150_io_hit; // @[cam.scala 93:27]
  wire  _io_hit_T_179 = _io_hit_T_149 | CAMLine_151_io_hit | CAMLine_152_io_hit | CAMLine_153_io_hit |
    CAMLine_154_io_hit | CAMLine_155_io_hit | CAMLine_156_io_hit | CAMLine_157_io_hit | CAMLine_158_io_hit |
    CAMLine_159_io_hit | CAMLine_160_io_hit | CAMLine_161_io_hit | CAMLine_162_io_hit | CAMLine_163_io_hit |
    CAMLine_164_io_hit | CAMLine_165_io_hit | CAMLine_166_io_hit | CAMLine_167_io_hit | CAMLine_168_io_hit |
    CAMLine_169_io_hit | CAMLine_170_io_hit | CAMLine_171_io_hit | CAMLine_172_io_hit | CAMLine_173_io_hit |
    CAMLine_174_io_hit | CAMLine_175_io_hit | CAMLine_176_io_hit | CAMLine_177_io_hit | CAMLine_178_io_hit |
    CAMLine_179_io_hit | CAMLine_180_io_hit; // @[cam.scala 93:27]
  wire  _io_hit_T_209 = _io_hit_T_179 | CAMLine_181_io_hit | CAMLine_182_io_hit | CAMLine_183_io_hit |
    CAMLine_184_io_hit | CAMLine_185_io_hit | CAMLine_186_io_hit | CAMLine_187_io_hit | CAMLine_188_io_hit |
    CAMLine_189_io_hit | CAMLine_190_io_hit | CAMLine_191_io_hit | CAMLine_192_io_hit | CAMLine_193_io_hit |
    CAMLine_194_io_hit | CAMLine_195_io_hit | CAMLine_196_io_hit | CAMLine_197_io_hit | CAMLine_198_io_hit |
    CAMLine_199_io_hit | CAMLine_200_io_hit | CAMLine_201_io_hit | CAMLine_202_io_hit | CAMLine_203_io_hit |
    CAMLine_204_io_hit | CAMLine_205_io_hit | CAMLine_206_io_hit | CAMLine_207_io_hit | CAMLine_208_io_hit |
    CAMLine_209_io_hit | CAMLine_210_io_hit; // @[cam.scala 93:27]
  wire  _io_hit_T_239 = _io_hit_T_209 | CAMLine_211_io_hit | CAMLine_212_io_hit | CAMLine_213_io_hit |
    CAMLine_214_io_hit | CAMLine_215_io_hit | CAMLine_216_io_hit | CAMLine_217_io_hit | CAMLine_218_io_hit |
    CAMLine_219_io_hit | CAMLine_220_io_hit | CAMLine_221_io_hit | CAMLine_222_io_hit | CAMLine_223_io_hit |
    CAMLine_224_io_hit | CAMLine_225_io_hit | CAMLine_226_io_hit | CAMLine_227_io_hit | CAMLine_228_io_hit |
    CAMLine_229_io_hit | CAMLine_230_io_hit | CAMLine_231_io_hit | CAMLine_232_io_hit | CAMLine_233_io_hit |
    CAMLine_234_io_hit | CAMLine_235_io_hit | CAMLine_236_io_hit | CAMLine_237_io_hit | CAMLine_238_io_hit |
    CAMLine_239_io_hit | CAMLine_240_io_hit; // @[cam.scala 93:27]
  CAMLine CAMLine ( // @[cam.scala 81:36]
    .clock(CAMLine_clock),
    .io_we(CAMLine_io_we),
    .io_wi(CAMLine_io_wi),
    .io_key(CAMLine_io_key),
    .io_din(CAMLine_io_din),
    .io_hit(CAMLine_io_hit)
  );
  CAMLine CAMLine_1 ( // @[cam.scala 81:36]
    .clock(CAMLine_1_clock),
    .io_we(CAMLine_1_io_we),
    .io_wi(CAMLine_1_io_wi),
    .io_key(CAMLine_1_io_key),
    .io_din(CAMLine_1_io_din),
    .io_hit(CAMLine_1_io_hit)
  );
  CAMLine CAMLine_2 ( // @[cam.scala 81:36]
    .clock(CAMLine_2_clock),
    .io_we(CAMLine_2_io_we),
    .io_wi(CAMLine_2_io_wi),
    .io_key(CAMLine_2_io_key),
    .io_din(CAMLine_2_io_din),
    .io_hit(CAMLine_2_io_hit)
  );
  CAMLine CAMLine_3 ( // @[cam.scala 81:36]
    .clock(CAMLine_3_clock),
    .io_we(CAMLine_3_io_we),
    .io_wi(CAMLine_3_io_wi),
    .io_key(CAMLine_3_io_key),
    .io_din(CAMLine_3_io_din),
    .io_hit(CAMLine_3_io_hit)
  );
  CAMLine CAMLine_4 ( // @[cam.scala 81:36]
    .clock(CAMLine_4_clock),
    .io_we(CAMLine_4_io_we),
    .io_wi(CAMLine_4_io_wi),
    .io_key(CAMLine_4_io_key),
    .io_din(CAMLine_4_io_din),
    .io_hit(CAMLine_4_io_hit)
  );
  CAMLine CAMLine_5 ( // @[cam.scala 81:36]
    .clock(CAMLine_5_clock),
    .io_we(CAMLine_5_io_we),
    .io_wi(CAMLine_5_io_wi),
    .io_key(CAMLine_5_io_key),
    .io_din(CAMLine_5_io_din),
    .io_hit(CAMLine_5_io_hit)
  );
  CAMLine CAMLine_6 ( // @[cam.scala 81:36]
    .clock(CAMLine_6_clock),
    .io_we(CAMLine_6_io_we),
    .io_wi(CAMLine_6_io_wi),
    .io_key(CAMLine_6_io_key),
    .io_din(CAMLine_6_io_din),
    .io_hit(CAMLine_6_io_hit)
  );
  CAMLine CAMLine_7 ( // @[cam.scala 81:36]
    .clock(CAMLine_7_clock),
    .io_we(CAMLine_7_io_we),
    .io_wi(CAMLine_7_io_wi),
    .io_key(CAMLine_7_io_key),
    .io_din(CAMLine_7_io_din),
    .io_hit(CAMLine_7_io_hit)
  );
  CAMLine CAMLine_8 ( // @[cam.scala 81:36]
    .clock(CAMLine_8_clock),
    .io_we(CAMLine_8_io_we),
    .io_wi(CAMLine_8_io_wi),
    .io_key(CAMLine_8_io_key),
    .io_din(CAMLine_8_io_din),
    .io_hit(CAMLine_8_io_hit)
  );
  CAMLine CAMLine_9 ( // @[cam.scala 81:36]
    .clock(CAMLine_9_clock),
    .io_we(CAMLine_9_io_we),
    .io_wi(CAMLine_9_io_wi),
    .io_key(CAMLine_9_io_key),
    .io_din(CAMLine_9_io_din),
    .io_hit(CAMLine_9_io_hit)
  );
  CAMLine CAMLine_10 ( // @[cam.scala 81:36]
    .clock(CAMLine_10_clock),
    .io_we(CAMLine_10_io_we),
    .io_wi(CAMLine_10_io_wi),
    .io_key(CAMLine_10_io_key),
    .io_din(CAMLine_10_io_din),
    .io_hit(CAMLine_10_io_hit)
  );
  CAMLine CAMLine_11 ( // @[cam.scala 81:36]
    .clock(CAMLine_11_clock),
    .io_we(CAMLine_11_io_we),
    .io_wi(CAMLine_11_io_wi),
    .io_key(CAMLine_11_io_key),
    .io_din(CAMLine_11_io_din),
    .io_hit(CAMLine_11_io_hit)
  );
  CAMLine CAMLine_12 ( // @[cam.scala 81:36]
    .clock(CAMLine_12_clock),
    .io_we(CAMLine_12_io_we),
    .io_wi(CAMLine_12_io_wi),
    .io_key(CAMLine_12_io_key),
    .io_din(CAMLine_12_io_din),
    .io_hit(CAMLine_12_io_hit)
  );
  CAMLine CAMLine_13 ( // @[cam.scala 81:36]
    .clock(CAMLine_13_clock),
    .io_we(CAMLine_13_io_we),
    .io_wi(CAMLine_13_io_wi),
    .io_key(CAMLine_13_io_key),
    .io_din(CAMLine_13_io_din),
    .io_hit(CAMLine_13_io_hit)
  );
  CAMLine CAMLine_14 ( // @[cam.scala 81:36]
    .clock(CAMLine_14_clock),
    .io_we(CAMLine_14_io_we),
    .io_wi(CAMLine_14_io_wi),
    .io_key(CAMLine_14_io_key),
    .io_din(CAMLine_14_io_din),
    .io_hit(CAMLine_14_io_hit)
  );
  CAMLine CAMLine_15 ( // @[cam.scala 81:36]
    .clock(CAMLine_15_clock),
    .io_we(CAMLine_15_io_we),
    .io_wi(CAMLine_15_io_wi),
    .io_key(CAMLine_15_io_key),
    .io_din(CAMLine_15_io_din),
    .io_hit(CAMLine_15_io_hit)
  );
  CAMLine CAMLine_16 ( // @[cam.scala 81:36]
    .clock(CAMLine_16_clock),
    .io_we(CAMLine_16_io_we),
    .io_wi(CAMLine_16_io_wi),
    .io_key(CAMLine_16_io_key),
    .io_din(CAMLine_16_io_din),
    .io_hit(CAMLine_16_io_hit)
  );
  CAMLine CAMLine_17 ( // @[cam.scala 81:36]
    .clock(CAMLine_17_clock),
    .io_we(CAMLine_17_io_we),
    .io_wi(CAMLine_17_io_wi),
    .io_key(CAMLine_17_io_key),
    .io_din(CAMLine_17_io_din),
    .io_hit(CAMLine_17_io_hit)
  );
  CAMLine CAMLine_18 ( // @[cam.scala 81:36]
    .clock(CAMLine_18_clock),
    .io_we(CAMLine_18_io_we),
    .io_wi(CAMLine_18_io_wi),
    .io_key(CAMLine_18_io_key),
    .io_din(CAMLine_18_io_din),
    .io_hit(CAMLine_18_io_hit)
  );
  CAMLine CAMLine_19 ( // @[cam.scala 81:36]
    .clock(CAMLine_19_clock),
    .io_we(CAMLine_19_io_we),
    .io_wi(CAMLine_19_io_wi),
    .io_key(CAMLine_19_io_key),
    .io_din(CAMLine_19_io_din),
    .io_hit(CAMLine_19_io_hit)
  );
  CAMLine CAMLine_20 ( // @[cam.scala 81:36]
    .clock(CAMLine_20_clock),
    .io_we(CAMLine_20_io_we),
    .io_wi(CAMLine_20_io_wi),
    .io_key(CAMLine_20_io_key),
    .io_din(CAMLine_20_io_din),
    .io_hit(CAMLine_20_io_hit)
  );
  CAMLine CAMLine_21 ( // @[cam.scala 81:36]
    .clock(CAMLine_21_clock),
    .io_we(CAMLine_21_io_we),
    .io_wi(CAMLine_21_io_wi),
    .io_key(CAMLine_21_io_key),
    .io_din(CAMLine_21_io_din),
    .io_hit(CAMLine_21_io_hit)
  );
  CAMLine CAMLine_22 ( // @[cam.scala 81:36]
    .clock(CAMLine_22_clock),
    .io_we(CAMLine_22_io_we),
    .io_wi(CAMLine_22_io_wi),
    .io_key(CAMLine_22_io_key),
    .io_din(CAMLine_22_io_din),
    .io_hit(CAMLine_22_io_hit)
  );
  CAMLine CAMLine_23 ( // @[cam.scala 81:36]
    .clock(CAMLine_23_clock),
    .io_we(CAMLine_23_io_we),
    .io_wi(CAMLine_23_io_wi),
    .io_key(CAMLine_23_io_key),
    .io_din(CAMLine_23_io_din),
    .io_hit(CAMLine_23_io_hit)
  );
  CAMLine CAMLine_24 ( // @[cam.scala 81:36]
    .clock(CAMLine_24_clock),
    .io_we(CAMLine_24_io_we),
    .io_wi(CAMLine_24_io_wi),
    .io_key(CAMLine_24_io_key),
    .io_din(CAMLine_24_io_din),
    .io_hit(CAMLine_24_io_hit)
  );
  CAMLine CAMLine_25 ( // @[cam.scala 81:36]
    .clock(CAMLine_25_clock),
    .io_we(CAMLine_25_io_we),
    .io_wi(CAMLine_25_io_wi),
    .io_key(CAMLine_25_io_key),
    .io_din(CAMLine_25_io_din),
    .io_hit(CAMLine_25_io_hit)
  );
  CAMLine CAMLine_26 ( // @[cam.scala 81:36]
    .clock(CAMLine_26_clock),
    .io_we(CAMLine_26_io_we),
    .io_wi(CAMLine_26_io_wi),
    .io_key(CAMLine_26_io_key),
    .io_din(CAMLine_26_io_din),
    .io_hit(CAMLine_26_io_hit)
  );
  CAMLine CAMLine_27 ( // @[cam.scala 81:36]
    .clock(CAMLine_27_clock),
    .io_we(CAMLine_27_io_we),
    .io_wi(CAMLine_27_io_wi),
    .io_key(CAMLine_27_io_key),
    .io_din(CAMLine_27_io_din),
    .io_hit(CAMLine_27_io_hit)
  );
  CAMLine CAMLine_28 ( // @[cam.scala 81:36]
    .clock(CAMLine_28_clock),
    .io_we(CAMLine_28_io_we),
    .io_wi(CAMLine_28_io_wi),
    .io_key(CAMLine_28_io_key),
    .io_din(CAMLine_28_io_din),
    .io_hit(CAMLine_28_io_hit)
  );
  CAMLine CAMLine_29 ( // @[cam.scala 81:36]
    .clock(CAMLine_29_clock),
    .io_we(CAMLine_29_io_we),
    .io_wi(CAMLine_29_io_wi),
    .io_key(CAMLine_29_io_key),
    .io_din(CAMLine_29_io_din),
    .io_hit(CAMLine_29_io_hit)
  );
  CAMLine CAMLine_30 ( // @[cam.scala 81:36]
    .clock(CAMLine_30_clock),
    .io_we(CAMLine_30_io_we),
    .io_wi(CAMLine_30_io_wi),
    .io_key(CAMLine_30_io_key),
    .io_din(CAMLine_30_io_din),
    .io_hit(CAMLine_30_io_hit)
  );
  CAMLine CAMLine_31 ( // @[cam.scala 81:36]
    .clock(CAMLine_31_clock),
    .io_we(CAMLine_31_io_we),
    .io_wi(CAMLine_31_io_wi),
    .io_key(CAMLine_31_io_key),
    .io_din(CAMLine_31_io_din),
    .io_hit(CAMLine_31_io_hit)
  );
  CAMLine CAMLine_32 ( // @[cam.scala 81:36]
    .clock(CAMLine_32_clock),
    .io_we(CAMLine_32_io_we),
    .io_wi(CAMLine_32_io_wi),
    .io_key(CAMLine_32_io_key),
    .io_din(CAMLine_32_io_din),
    .io_hit(CAMLine_32_io_hit)
  );
  CAMLine CAMLine_33 ( // @[cam.scala 81:36]
    .clock(CAMLine_33_clock),
    .io_we(CAMLine_33_io_we),
    .io_wi(CAMLine_33_io_wi),
    .io_key(CAMLine_33_io_key),
    .io_din(CAMLine_33_io_din),
    .io_hit(CAMLine_33_io_hit)
  );
  CAMLine CAMLine_34 ( // @[cam.scala 81:36]
    .clock(CAMLine_34_clock),
    .io_we(CAMLine_34_io_we),
    .io_wi(CAMLine_34_io_wi),
    .io_key(CAMLine_34_io_key),
    .io_din(CAMLine_34_io_din),
    .io_hit(CAMLine_34_io_hit)
  );
  CAMLine CAMLine_35 ( // @[cam.scala 81:36]
    .clock(CAMLine_35_clock),
    .io_we(CAMLine_35_io_we),
    .io_wi(CAMLine_35_io_wi),
    .io_key(CAMLine_35_io_key),
    .io_din(CAMLine_35_io_din),
    .io_hit(CAMLine_35_io_hit)
  );
  CAMLine CAMLine_36 ( // @[cam.scala 81:36]
    .clock(CAMLine_36_clock),
    .io_we(CAMLine_36_io_we),
    .io_wi(CAMLine_36_io_wi),
    .io_key(CAMLine_36_io_key),
    .io_din(CAMLine_36_io_din),
    .io_hit(CAMLine_36_io_hit)
  );
  CAMLine CAMLine_37 ( // @[cam.scala 81:36]
    .clock(CAMLine_37_clock),
    .io_we(CAMLine_37_io_we),
    .io_wi(CAMLine_37_io_wi),
    .io_key(CAMLine_37_io_key),
    .io_din(CAMLine_37_io_din),
    .io_hit(CAMLine_37_io_hit)
  );
  CAMLine CAMLine_38 ( // @[cam.scala 81:36]
    .clock(CAMLine_38_clock),
    .io_we(CAMLine_38_io_we),
    .io_wi(CAMLine_38_io_wi),
    .io_key(CAMLine_38_io_key),
    .io_din(CAMLine_38_io_din),
    .io_hit(CAMLine_38_io_hit)
  );
  CAMLine CAMLine_39 ( // @[cam.scala 81:36]
    .clock(CAMLine_39_clock),
    .io_we(CAMLine_39_io_we),
    .io_wi(CAMLine_39_io_wi),
    .io_key(CAMLine_39_io_key),
    .io_din(CAMLine_39_io_din),
    .io_hit(CAMLine_39_io_hit)
  );
  CAMLine CAMLine_40 ( // @[cam.scala 81:36]
    .clock(CAMLine_40_clock),
    .io_we(CAMLine_40_io_we),
    .io_wi(CAMLine_40_io_wi),
    .io_key(CAMLine_40_io_key),
    .io_din(CAMLine_40_io_din),
    .io_hit(CAMLine_40_io_hit)
  );
  CAMLine CAMLine_41 ( // @[cam.scala 81:36]
    .clock(CAMLine_41_clock),
    .io_we(CAMLine_41_io_we),
    .io_wi(CAMLine_41_io_wi),
    .io_key(CAMLine_41_io_key),
    .io_din(CAMLine_41_io_din),
    .io_hit(CAMLine_41_io_hit)
  );
  CAMLine CAMLine_42 ( // @[cam.scala 81:36]
    .clock(CAMLine_42_clock),
    .io_we(CAMLine_42_io_we),
    .io_wi(CAMLine_42_io_wi),
    .io_key(CAMLine_42_io_key),
    .io_din(CAMLine_42_io_din),
    .io_hit(CAMLine_42_io_hit)
  );
  CAMLine CAMLine_43 ( // @[cam.scala 81:36]
    .clock(CAMLine_43_clock),
    .io_we(CAMLine_43_io_we),
    .io_wi(CAMLine_43_io_wi),
    .io_key(CAMLine_43_io_key),
    .io_din(CAMLine_43_io_din),
    .io_hit(CAMLine_43_io_hit)
  );
  CAMLine CAMLine_44 ( // @[cam.scala 81:36]
    .clock(CAMLine_44_clock),
    .io_we(CAMLine_44_io_we),
    .io_wi(CAMLine_44_io_wi),
    .io_key(CAMLine_44_io_key),
    .io_din(CAMLine_44_io_din),
    .io_hit(CAMLine_44_io_hit)
  );
  CAMLine CAMLine_45 ( // @[cam.scala 81:36]
    .clock(CAMLine_45_clock),
    .io_we(CAMLine_45_io_we),
    .io_wi(CAMLine_45_io_wi),
    .io_key(CAMLine_45_io_key),
    .io_din(CAMLine_45_io_din),
    .io_hit(CAMLine_45_io_hit)
  );
  CAMLine CAMLine_46 ( // @[cam.scala 81:36]
    .clock(CAMLine_46_clock),
    .io_we(CAMLine_46_io_we),
    .io_wi(CAMLine_46_io_wi),
    .io_key(CAMLine_46_io_key),
    .io_din(CAMLine_46_io_din),
    .io_hit(CAMLine_46_io_hit)
  );
  CAMLine CAMLine_47 ( // @[cam.scala 81:36]
    .clock(CAMLine_47_clock),
    .io_we(CAMLine_47_io_we),
    .io_wi(CAMLine_47_io_wi),
    .io_key(CAMLine_47_io_key),
    .io_din(CAMLine_47_io_din),
    .io_hit(CAMLine_47_io_hit)
  );
  CAMLine CAMLine_48 ( // @[cam.scala 81:36]
    .clock(CAMLine_48_clock),
    .io_we(CAMLine_48_io_we),
    .io_wi(CAMLine_48_io_wi),
    .io_key(CAMLine_48_io_key),
    .io_din(CAMLine_48_io_din),
    .io_hit(CAMLine_48_io_hit)
  );
  CAMLine CAMLine_49 ( // @[cam.scala 81:36]
    .clock(CAMLine_49_clock),
    .io_we(CAMLine_49_io_we),
    .io_wi(CAMLine_49_io_wi),
    .io_key(CAMLine_49_io_key),
    .io_din(CAMLine_49_io_din),
    .io_hit(CAMLine_49_io_hit)
  );
  CAMLine CAMLine_50 ( // @[cam.scala 81:36]
    .clock(CAMLine_50_clock),
    .io_we(CAMLine_50_io_we),
    .io_wi(CAMLine_50_io_wi),
    .io_key(CAMLine_50_io_key),
    .io_din(CAMLine_50_io_din),
    .io_hit(CAMLine_50_io_hit)
  );
  CAMLine CAMLine_51 ( // @[cam.scala 81:36]
    .clock(CAMLine_51_clock),
    .io_we(CAMLine_51_io_we),
    .io_wi(CAMLine_51_io_wi),
    .io_key(CAMLine_51_io_key),
    .io_din(CAMLine_51_io_din),
    .io_hit(CAMLine_51_io_hit)
  );
  CAMLine CAMLine_52 ( // @[cam.scala 81:36]
    .clock(CAMLine_52_clock),
    .io_we(CAMLine_52_io_we),
    .io_wi(CAMLine_52_io_wi),
    .io_key(CAMLine_52_io_key),
    .io_din(CAMLine_52_io_din),
    .io_hit(CAMLine_52_io_hit)
  );
  CAMLine CAMLine_53 ( // @[cam.scala 81:36]
    .clock(CAMLine_53_clock),
    .io_we(CAMLine_53_io_we),
    .io_wi(CAMLine_53_io_wi),
    .io_key(CAMLine_53_io_key),
    .io_din(CAMLine_53_io_din),
    .io_hit(CAMLine_53_io_hit)
  );
  CAMLine CAMLine_54 ( // @[cam.scala 81:36]
    .clock(CAMLine_54_clock),
    .io_we(CAMLine_54_io_we),
    .io_wi(CAMLine_54_io_wi),
    .io_key(CAMLine_54_io_key),
    .io_din(CAMLine_54_io_din),
    .io_hit(CAMLine_54_io_hit)
  );
  CAMLine CAMLine_55 ( // @[cam.scala 81:36]
    .clock(CAMLine_55_clock),
    .io_we(CAMLine_55_io_we),
    .io_wi(CAMLine_55_io_wi),
    .io_key(CAMLine_55_io_key),
    .io_din(CAMLine_55_io_din),
    .io_hit(CAMLine_55_io_hit)
  );
  CAMLine CAMLine_56 ( // @[cam.scala 81:36]
    .clock(CAMLine_56_clock),
    .io_we(CAMLine_56_io_we),
    .io_wi(CAMLine_56_io_wi),
    .io_key(CAMLine_56_io_key),
    .io_din(CAMLine_56_io_din),
    .io_hit(CAMLine_56_io_hit)
  );
  CAMLine CAMLine_57 ( // @[cam.scala 81:36]
    .clock(CAMLine_57_clock),
    .io_we(CAMLine_57_io_we),
    .io_wi(CAMLine_57_io_wi),
    .io_key(CAMLine_57_io_key),
    .io_din(CAMLine_57_io_din),
    .io_hit(CAMLine_57_io_hit)
  );
  CAMLine CAMLine_58 ( // @[cam.scala 81:36]
    .clock(CAMLine_58_clock),
    .io_we(CAMLine_58_io_we),
    .io_wi(CAMLine_58_io_wi),
    .io_key(CAMLine_58_io_key),
    .io_din(CAMLine_58_io_din),
    .io_hit(CAMLine_58_io_hit)
  );
  CAMLine CAMLine_59 ( // @[cam.scala 81:36]
    .clock(CAMLine_59_clock),
    .io_we(CAMLine_59_io_we),
    .io_wi(CAMLine_59_io_wi),
    .io_key(CAMLine_59_io_key),
    .io_din(CAMLine_59_io_din),
    .io_hit(CAMLine_59_io_hit)
  );
  CAMLine CAMLine_60 ( // @[cam.scala 81:36]
    .clock(CAMLine_60_clock),
    .io_we(CAMLine_60_io_we),
    .io_wi(CAMLine_60_io_wi),
    .io_key(CAMLine_60_io_key),
    .io_din(CAMLine_60_io_din),
    .io_hit(CAMLine_60_io_hit)
  );
  CAMLine CAMLine_61 ( // @[cam.scala 81:36]
    .clock(CAMLine_61_clock),
    .io_we(CAMLine_61_io_we),
    .io_wi(CAMLine_61_io_wi),
    .io_key(CAMLine_61_io_key),
    .io_din(CAMLine_61_io_din),
    .io_hit(CAMLine_61_io_hit)
  );
  CAMLine CAMLine_62 ( // @[cam.scala 81:36]
    .clock(CAMLine_62_clock),
    .io_we(CAMLine_62_io_we),
    .io_wi(CAMLine_62_io_wi),
    .io_key(CAMLine_62_io_key),
    .io_din(CAMLine_62_io_din),
    .io_hit(CAMLine_62_io_hit)
  );
  CAMLine CAMLine_63 ( // @[cam.scala 81:36]
    .clock(CAMLine_63_clock),
    .io_we(CAMLine_63_io_we),
    .io_wi(CAMLine_63_io_wi),
    .io_key(CAMLine_63_io_key),
    .io_din(CAMLine_63_io_din),
    .io_hit(CAMLine_63_io_hit)
  );
  CAMLine CAMLine_64 ( // @[cam.scala 81:36]
    .clock(CAMLine_64_clock),
    .io_we(CAMLine_64_io_we),
    .io_wi(CAMLine_64_io_wi),
    .io_key(CAMLine_64_io_key),
    .io_din(CAMLine_64_io_din),
    .io_hit(CAMLine_64_io_hit)
  );
  CAMLine CAMLine_65 ( // @[cam.scala 81:36]
    .clock(CAMLine_65_clock),
    .io_we(CAMLine_65_io_we),
    .io_wi(CAMLine_65_io_wi),
    .io_key(CAMLine_65_io_key),
    .io_din(CAMLine_65_io_din),
    .io_hit(CAMLine_65_io_hit)
  );
  CAMLine CAMLine_66 ( // @[cam.scala 81:36]
    .clock(CAMLine_66_clock),
    .io_we(CAMLine_66_io_we),
    .io_wi(CAMLine_66_io_wi),
    .io_key(CAMLine_66_io_key),
    .io_din(CAMLine_66_io_din),
    .io_hit(CAMLine_66_io_hit)
  );
  CAMLine CAMLine_67 ( // @[cam.scala 81:36]
    .clock(CAMLine_67_clock),
    .io_we(CAMLine_67_io_we),
    .io_wi(CAMLine_67_io_wi),
    .io_key(CAMLine_67_io_key),
    .io_din(CAMLine_67_io_din),
    .io_hit(CAMLine_67_io_hit)
  );
  CAMLine CAMLine_68 ( // @[cam.scala 81:36]
    .clock(CAMLine_68_clock),
    .io_we(CAMLine_68_io_we),
    .io_wi(CAMLine_68_io_wi),
    .io_key(CAMLine_68_io_key),
    .io_din(CAMLine_68_io_din),
    .io_hit(CAMLine_68_io_hit)
  );
  CAMLine CAMLine_69 ( // @[cam.scala 81:36]
    .clock(CAMLine_69_clock),
    .io_we(CAMLine_69_io_we),
    .io_wi(CAMLine_69_io_wi),
    .io_key(CAMLine_69_io_key),
    .io_din(CAMLine_69_io_din),
    .io_hit(CAMLine_69_io_hit)
  );
  CAMLine CAMLine_70 ( // @[cam.scala 81:36]
    .clock(CAMLine_70_clock),
    .io_we(CAMLine_70_io_we),
    .io_wi(CAMLine_70_io_wi),
    .io_key(CAMLine_70_io_key),
    .io_din(CAMLine_70_io_din),
    .io_hit(CAMLine_70_io_hit)
  );
  CAMLine CAMLine_71 ( // @[cam.scala 81:36]
    .clock(CAMLine_71_clock),
    .io_we(CAMLine_71_io_we),
    .io_wi(CAMLine_71_io_wi),
    .io_key(CAMLine_71_io_key),
    .io_din(CAMLine_71_io_din),
    .io_hit(CAMLine_71_io_hit)
  );
  CAMLine CAMLine_72 ( // @[cam.scala 81:36]
    .clock(CAMLine_72_clock),
    .io_we(CAMLine_72_io_we),
    .io_wi(CAMLine_72_io_wi),
    .io_key(CAMLine_72_io_key),
    .io_din(CAMLine_72_io_din),
    .io_hit(CAMLine_72_io_hit)
  );
  CAMLine CAMLine_73 ( // @[cam.scala 81:36]
    .clock(CAMLine_73_clock),
    .io_we(CAMLine_73_io_we),
    .io_wi(CAMLine_73_io_wi),
    .io_key(CAMLine_73_io_key),
    .io_din(CAMLine_73_io_din),
    .io_hit(CAMLine_73_io_hit)
  );
  CAMLine CAMLine_74 ( // @[cam.scala 81:36]
    .clock(CAMLine_74_clock),
    .io_we(CAMLine_74_io_we),
    .io_wi(CAMLine_74_io_wi),
    .io_key(CAMLine_74_io_key),
    .io_din(CAMLine_74_io_din),
    .io_hit(CAMLine_74_io_hit)
  );
  CAMLine CAMLine_75 ( // @[cam.scala 81:36]
    .clock(CAMLine_75_clock),
    .io_we(CAMLine_75_io_we),
    .io_wi(CAMLine_75_io_wi),
    .io_key(CAMLine_75_io_key),
    .io_din(CAMLine_75_io_din),
    .io_hit(CAMLine_75_io_hit)
  );
  CAMLine CAMLine_76 ( // @[cam.scala 81:36]
    .clock(CAMLine_76_clock),
    .io_we(CAMLine_76_io_we),
    .io_wi(CAMLine_76_io_wi),
    .io_key(CAMLine_76_io_key),
    .io_din(CAMLine_76_io_din),
    .io_hit(CAMLine_76_io_hit)
  );
  CAMLine CAMLine_77 ( // @[cam.scala 81:36]
    .clock(CAMLine_77_clock),
    .io_we(CAMLine_77_io_we),
    .io_wi(CAMLine_77_io_wi),
    .io_key(CAMLine_77_io_key),
    .io_din(CAMLine_77_io_din),
    .io_hit(CAMLine_77_io_hit)
  );
  CAMLine CAMLine_78 ( // @[cam.scala 81:36]
    .clock(CAMLine_78_clock),
    .io_we(CAMLine_78_io_we),
    .io_wi(CAMLine_78_io_wi),
    .io_key(CAMLine_78_io_key),
    .io_din(CAMLine_78_io_din),
    .io_hit(CAMLine_78_io_hit)
  );
  CAMLine CAMLine_79 ( // @[cam.scala 81:36]
    .clock(CAMLine_79_clock),
    .io_we(CAMLine_79_io_we),
    .io_wi(CAMLine_79_io_wi),
    .io_key(CAMLine_79_io_key),
    .io_din(CAMLine_79_io_din),
    .io_hit(CAMLine_79_io_hit)
  );
  CAMLine CAMLine_80 ( // @[cam.scala 81:36]
    .clock(CAMLine_80_clock),
    .io_we(CAMLine_80_io_we),
    .io_wi(CAMLine_80_io_wi),
    .io_key(CAMLine_80_io_key),
    .io_din(CAMLine_80_io_din),
    .io_hit(CAMLine_80_io_hit)
  );
  CAMLine CAMLine_81 ( // @[cam.scala 81:36]
    .clock(CAMLine_81_clock),
    .io_we(CAMLine_81_io_we),
    .io_wi(CAMLine_81_io_wi),
    .io_key(CAMLine_81_io_key),
    .io_din(CAMLine_81_io_din),
    .io_hit(CAMLine_81_io_hit)
  );
  CAMLine CAMLine_82 ( // @[cam.scala 81:36]
    .clock(CAMLine_82_clock),
    .io_we(CAMLine_82_io_we),
    .io_wi(CAMLine_82_io_wi),
    .io_key(CAMLine_82_io_key),
    .io_din(CAMLine_82_io_din),
    .io_hit(CAMLine_82_io_hit)
  );
  CAMLine CAMLine_83 ( // @[cam.scala 81:36]
    .clock(CAMLine_83_clock),
    .io_we(CAMLine_83_io_we),
    .io_wi(CAMLine_83_io_wi),
    .io_key(CAMLine_83_io_key),
    .io_din(CAMLine_83_io_din),
    .io_hit(CAMLine_83_io_hit)
  );
  CAMLine CAMLine_84 ( // @[cam.scala 81:36]
    .clock(CAMLine_84_clock),
    .io_we(CAMLine_84_io_we),
    .io_wi(CAMLine_84_io_wi),
    .io_key(CAMLine_84_io_key),
    .io_din(CAMLine_84_io_din),
    .io_hit(CAMLine_84_io_hit)
  );
  CAMLine CAMLine_85 ( // @[cam.scala 81:36]
    .clock(CAMLine_85_clock),
    .io_we(CAMLine_85_io_we),
    .io_wi(CAMLine_85_io_wi),
    .io_key(CAMLine_85_io_key),
    .io_din(CAMLine_85_io_din),
    .io_hit(CAMLine_85_io_hit)
  );
  CAMLine CAMLine_86 ( // @[cam.scala 81:36]
    .clock(CAMLine_86_clock),
    .io_we(CAMLine_86_io_we),
    .io_wi(CAMLine_86_io_wi),
    .io_key(CAMLine_86_io_key),
    .io_din(CAMLine_86_io_din),
    .io_hit(CAMLine_86_io_hit)
  );
  CAMLine CAMLine_87 ( // @[cam.scala 81:36]
    .clock(CAMLine_87_clock),
    .io_we(CAMLine_87_io_we),
    .io_wi(CAMLine_87_io_wi),
    .io_key(CAMLine_87_io_key),
    .io_din(CAMLine_87_io_din),
    .io_hit(CAMLine_87_io_hit)
  );
  CAMLine CAMLine_88 ( // @[cam.scala 81:36]
    .clock(CAMLine_88_clock),
    .io_we(CAMLine_88_io_we),
    .io_wi(CAMLine_88_io_wi),
    .io_key(CAMLine_88_io_key),
    .io_din(CAMLine_88_io_din),
    .io_hit(CAMLine_88_io_hit)
  );
  CAMLine CAMLine_89 ( // @[cam.scala 81:36]
    .clock(CAMLine_89_clock),
    .io_we(CAMLine_89_io_we),
    .io_wi(CAMLine_89_io_wi),
    .io_key(CAMLine_89_io_key),
    .io_din(CAMLine_89_io_din),
    .io_hit(CAMLine_89_io_hit)
  );
  CAMLine CAMLine_90 ( // @[cam.scala 81:36]
    .clock(CAMLine_90_clock),
    .io_we(CAMLine_90_io_we),
    .io_wi(CAMLine_90_io_wi),
    .io_key(CAMLine_90_io_key),
    .io_din(CAMLine_90_io_din),
    .io_hit(CAMLine_90_io_hit)
  );
  CAMLine CAMLine_91 ( // @[cam.scala 81:36]
    .clock(CAMLine_91_clock),
    .io_we(CAMLine_91_io_we),
    .io_wi(CAMLine_91_io_wi),
    .io_key(CAMLine_91_io_key),
    .io_din(CAMLine_91_io_din),
    .io_hit(CAMLine_91_io_hit)
  );
  CAMLine CAMLine_92 ( // @[cam.scala 81:36]
    .clock(CAMLine_92_clock),
    .io_we(CAMLine_92_io_we),
    .io_wi(CAMLine_92_io_wi),
    .io_key(CAMLine_92_io_key),
    .io_din(CAMLine_92_io_din),
    .io_hit(CAMLine_92_io_hit)
  );
  CAMLine CAMLine_93 ( // @[cam.scala 81:36]
    .clock(CAMLine_93_clock),
    .io_we(CAMLine_93_io_we),
    .io_wi(CAMLine_93_io_wi),
    .io_key(CAMLine_93_io_key),
    .io_din(CAMLine_93_io_din),
    .io_hit(CAMLine_93_io_hit)
  );
  CAMLine CAMLine_94 ( // @[cam.scala 81:36]
    .clock(CAMLine_94_clock),
    .io_we(CAMLine_94_io_we),
    .io_wi(CAMLine_94_io_wi),
    .io_key(CAMLine_94_io_key),
    .io_din(CAMLine_94_io_din),
    .io_hit(CAMLine_94_io_hit)
  );
  CAMLine CAMLine_95 ( // @[cam.scala 81:36]
    .clock(CAMLine_95_clock),
    .io_we(CAMLine_95_io_we),
    .io_wi(CAMLine_95_io_wi),
    .io_key(CAMLine_95_io_key),
    .io_din(CAMLine_95_io_din),
    .io_hit(CAMLine_95_io_hit)
  );
  CAMLine CAMLine_96 ( // @[cam.scala 81:36]
    .clock(CAMLine_96_clock),
    .io_we(CAMLine_96_io_we),
    .io_wi(CAMLine_96_io_wi),
    .io_key(CAMLine_96_io_key),
    .io_din(CAMLine_96_io_din),
    .io_hit(CAMLine_96_io_hit)
  );
  CAMLine CAMLine_97 ( // @[cam.scala 81:36]
    .clock(CAMLine_97_clock),
    .io_we(CAMLine_97_io_we),
    .io_wi(CAMLine_97_io_wi),
    .io_key(CAMLine_97_io_key),
    .io_din(CAMLine_97_io_din),
    .io_hit(CAMLine_97_io_hit)
  );
  CAMLine CAMLine_98 ( // @[cam.scala 81:36]
    .clock(CAMLine_98_clock),
    .io_we(CAMLine_98_io_we),
    .io_wi(CAMLine_98_io_wi),
    .io_key(CAMLine_98_io_key),
    .io_din(CAMLine_98_io_din),
    .io_hit(CAMLine_98_io_hit)
  );
  CAMLine CAMLine_99 ( // @[cam.scala 81:36]
    .clock(CAMLine_99_clock),
    .io_we(CAMLine_99_io_we),
    .io_wi(CAMLine_99_io_wi),
    .io_key(CAMLine_99_io_key),
    .io_din(CAMLine_99_io_din),
    .io_hit(CAMLine_99_io_hit)
  );
  CAMLine CAMLine_100 ( // @[cam.scala 81:36]
    .clock(CAMLine_100_clock),
    .io_we(CAMLine_100_io_we),
    .io_wi(CAMLine_100_io_wi),
    .io_key(CAMLine_100_io_key),
    .io_din(CAMLine_100_io_din),
    .io_hit(CAMLine_100_io_hit)
  );
  CAMLine CAMLine_101 ( // @[cam.scala 81:36]
    .clock(CAMLine_101_clock),
    .io_we(CAMLine_101_io_we),
    .io_wi(CAMLine_101_io_wi),
    .io_key(CAMLine_101_io_key),
    .io_din(CAMLine_101_io_din),
    .io_hit(CAMLine_101_io_hit)
  );
  CAMLine CAMLine_102 ( // @[cam.scala 81:36]
    .clock(CAMLine_102_clock),
    .io_we(CAMLine_102_io_we),
    .io_wi(CAMLine_102_io_wi),
    .io_key(CAMLine_102_io_key),
    .io_din(CAMLine_102_io_din),
    .io_hit(CAMLine_102_io_hit)
  );
  CAMLine CAMLine_103 ( // @[cam.scala 81:36]
    .clock(CAMLine_103_clock),
    .io_we(CAMLine_103_io_we),
    .io_wi(CAMLine_103_io_wi),
    .io_key(CAMLine_103_io_key),
    .io_din(CAMLine_103_io_din),
    .io_hit(CAMLine_103_io_hit)
  );
  CAMLine CAMLine_104 ( // @[cam.scala 81:36]
    .clock(CAMLine_104_clock),
    .io_we(CAMLine_104_io_we),
    .io_wi(CAMLine_104_io_wi),
    .io_key(CAMLine_104_io_key),
    .io_din(CAMLine_104_io_din),
    .io_hit(CAMLine_104_io_hit)
  );
  CAMLine CAMLine_105 ( // @[cam.scala 81:36]
    .clock(CAMLine_105_clock),
    .io_we(CAMLine_105_io_we),
    .io_wi(CAMLine_105_io_wi),
    .io_key(CAMLine_105_io_key),
    .io_din(CAMLine_105_io_din),
    .io_hit(CAMLine_105_io_hit)
  );
  CAMLine CAMLine_106 ( // @[cam.scala 81:36]
    .clock(CAMLine_106_clock),
    .io_we(CAMLine_106_io_we),
    .io_wi(CAMLine_106_io_wi),
    .io_key(CAMLine_106_io_key),
    .io_din(CAMLine_106_io_din),
    .io_hit(CAMLine_106_io_hit)
  );
  CAMLine CAMLine_107 ( // @[cam.scala 81:36]
    .clock(CAMLine_107_clock),
    .io_we(CAMLine_107_io_we),
    .io_wi(CAMLine_107_io_wi),
    .io_key(CAMLine_107_io_key),
    .io_din(CAMLine_107_io_din),
    .io_hit(CAMLine_107_io_hit)
  );
  CAMLine CAMLine_108 ( // @[cam.scala 81:36]
    .clock(CAMLine_108_clock),
    .io_we(CAMLine_108_io_we),
    .io_wi(CAMLine_108_io_wi),
    .io_key(CAMLine_108_io_key),
    .io_din(CAMLine_108_io_din),
    .io_hit(CAMLine_108_io_hit)
  );
  CAMLine CAMLine_109 ( // @[cam.scala 81:36]
    .clock(CAMLine_109_clock),
    .io_we(CAMLine_109_io_we),
    .io_wi(CAMLine_109_io_wi),
    .io_key(CAMLine_109_io_key),
    .io_din(CAMLine_109_io_din),
    .io_hit(CAMLine_109_io_hit)
  );
  CAMLine CAMLine_110 ( // @[cam.scala 81:36]
    .clock(CAMLine_110_clock),
    .io_we(CAMLine_110_io_we),
    .io_wi(CAMLine_110_io_wi),
    .io_key(CAMLine_110_io_key),
    .io_din(CAMLine_110_io_din),
    .io_hit(CAMLine_110_io_hit)
  );
  CAMLine CAMLine_111 ( // @[cam.scala 81:36]
    .clock(CAMLine_111_clock),
    .io_we(CAMLine_111_io_we),
    .io_wi(CAMLine_111_io_wi),
    .io_key(CAMLine_111_io_key),
    .io_din(CAMLine_111_io_din),
    .io_hit(CAMLine_111_io_hit)
  );
  CAMLine CAMLine_112 ( // @[cam.scala 81:36]
    .clock(CAMLine_112_clock),
    .io_we(CAMLine_112_io_we),
    .io_wi(CAMLine_112_io_wi),
    .io_key(CAMLine_112_io_key),
    .io_din(CAMLine_112_io_din),
    .io_hit(CAMLine_112_io_hit)
  );
  CAMLine CAMLine_113 ( // @[cam.scala 81:36]
    .clock(CAMLine_113_clock),
    .io_we(CAMLine_113_io_we),
    .io_wi(CAMLine_113_io_wi),
    .io_key(CAMLine_113_io_key),
    .io_din(CAMLine_113_io_din),
    .io_hit(CAMLine_113_io_hit)
  );
  CAMLine CAMLine_114 ( // @[cam.scala 81:36]
    .clock(CAMLine_114_clock),
    .io_we(CAMLine_114_io_we),
    .io_wi(CAMLine_114_io_wi),
    .io_key(CAMLine_114_io_key),
    .io_din(CAMLine_114_io_din),
    .io_hit(CAMLine_114_io_hit)
  );
  CAMLine CAMLine_115 ( // @[cam.scala 81:36]
    .clock(CAMLine_115_clock),
    .io_we(CAMLine_115_io_we),
    .io_wi(CAMLine_115_io_wi),
    .io_key(CAMLine_115_io_key),
    .io_din(CAMLine_115_io_din),
    .io_hit(CAMLine_115_io_hit)
  );
  CAMLine CAMLine_116 ( // @[cam.scala 81:36]
    .clock(CAMLine_116_clock),
    .io_we(CAMLine_116_io_we),
    .io_wi(CAMLine_116_io_wi),
    .io_key(CAMLine_116_io_key),
    .io_din(CAMLine_116_io_din),
    .io_hit(CAMLine_116_io_hit)
  );
  CAMLine CAMLine_117 ( // @[cam.scala 81:36]
    .clock(CAMLine_117_clock),
    .io_we(CAMLine_117_io_we),
    .io_wi(CAMLine_117_io_wi),
    .io_key(CAMLine_117_io_key),
    .io_din(CAMLine_117_io_din),
    .io_hit(CAMLine_117_io_hit)
  );
  CAMLine CAMLine_118 ( // @[cam.scala 81:36]
    .clock(CAMLine_118_clock),
    .io_we(CAMLine_118_io_we),
    .io_wi(CAMLine_118_io_wi),
    .io_key(CAMLine_118_io_key),
    .io_din(CAMLine_118_io_din),
    .io_hit(CAMLine_118_io_hit)
  );
  CAMLine CAMLine_119 ( // @[cam.scala 81:36]
    .clock(CAMLine_119_clock),
    .io_we(CAMLine_119_io_we),
    .io_wi(CAMLine_119_io_wi),
    .io_key(CAMLine_119_io_key),
    .io_din(CAMLine_119_io_din),
    .io_hit(CAMLine_119_io_hit)
  );
  CAMLine CAMLine_120 ( // @[cam.scala 81:36]
    .clock(CAMLine_120_clock),
    .io_we(CAMLine_120_io_we),
    .io_wi(CAMLine_120_io_wi),
    .io_key(CAMLine_120_io_key),
    .io_din(CAMLine_120_io_din),
    .io_hit(CAMLine_120_io_hit)
  );
  CAMLine CAMLine_121 ( // @[cam.scala 81:36]
    .clock(CAMLine_121_clock),
    .io_we(CAMLine_121_io_we),
    .io_wi(CAMLine_121_io_wi),
    .io_key(CAMLine_121_io_key),
    .io_din(CAMLine_121_io_din),
    .io_hit(CAMLine_121_io_hit)
  );
  CAMLine CAMLine_122 ( // @[cam.scala 81:36]
    .clock(CAMLine_122_clock),
    .io_we(CAMLine_122_io_we),
    .io_wi(CAMLine_122_io_wi),
    .io_key(CAMLine_122_io_key),
    .io_din(CAMLine_122_io_din),
    .io_hit(CAMLine_122_io_hit)
  );
  CAMLine CAMLine_123 ( // @[cam.scala 81:36]
    .clock(CAMLine_123_clock),
    .io_we(CAMLine_123_io_we),
    .io_wi(CAMLine_123_io_wi),
    .io_key(CAMLine_123_io_key),
    .io_din(CAMLine_123_io_din),
    .io_hit(CAMLine_123_io_hit)
  );
  CAMLine CAMLine_124 ( // @[cam.scala 81:36]
    .clock(CAMLine_124_clock),
    .io_we(CAMLine_124_io_we),
    .io_wi(CAMLine_124_io_wi),
    .io_key(CAMLine_124_io_key),
    .io_din(CAMLine_124_io_din),
    .io_hit(CAMLine_124_io_hit)
  );
  CAMLine CAMLine_125 ( // @[cam.scala 81:36]
    .clock(CAMLine_125_clock),
    .io_we(CAMLine_125_io_we),
    .io_wi(CAMLine_125_io_wi),
    .io_key(CAMLine_125_io_key),
    .io_din(CAMLine_125_io_din),
    .io_hit(CAMLine_125_io_hit)
  );
  CAMLine CAMLine_126 ( // @[cam.scala 81:36]
    .clock(CAMLine_126_clock),
    .io_we(CAMLine_126_io_we),
    .io_wi(CAMLine_126_io_wi),
    .io_key(CAMLine_126_io_key),
    .io_din(CAMLine_126_io_din),
    .io_hit(CAMLine_126_io_hit)
  );
  CAMLine CAMLine_127 ( // @[cam.scala 81:36]
    .clock(CAMLine_127_clock),
    .io_we(CAMLine_127_io_we),
    .io_wi(CAMLine_127_io_wi),
    .io_key(CAMLine_127_io_key),
    .io_din(CAMLine_127_io_din),
    .io_hit(CAMLine_127_io_hit)
  );
  CAMLine CAMLine_128 ( // @[cam.scala 81:36]
    .clock(CAMLine_128_clock),
    .io_we(CAMLine_128_io_we),
    .io_wi(CAMLine_128_io_wi),
    .io_key(CAMLine_128_io_key),
    .io_din(CAMLine_128_io_din),
    .io_hit(CAMLine_128_io_hit)
  );
  CAMLine CAMLine_129 ( // @[cam.scala 81:36]
    .clock(CAMLine_129_clock),
    .io_we(CAMLine_129_io_we),
    .io_wi(CAMLine_129_io_wi),
    .io_key(CAMLine_129_io_key),
    .io_din(CAMLine_129_io_din),
    .io_hit(CAMLine_129_io_hit)
  );
  CAMLine CAMLine_130 ( // @[cam.scala 81:36]
    .clock(CAMLine_130_clock),
    .io_we(CAMLine_130_io_we),
    .io_wi(CAMLine_130_io_wi),
    .io_key(CAMLine_130_io_key),
    .io_din(CAMLine_130_io_din),
    .io_hit(CAMLine_130_io_hit)
  );
  CAMLine CAMLine_131 ( // @[cam.scala 81:36]
    .clock(CAMLine_131_clock),
    .io_we(CAMLine_131_io_we),
    .io_wi(CAMLine_131_io_wi),
    .io_key(CAMLine_131_io_key),
    .io_din(CAMLine_131_io_din),
    .io_hit(CAMLine_131_io_hit)
  );
  CAMLine CAMLine_132 ( // @[cam.scala 81:36]
    .clock(CAMLine_132_clock),
    .io_we(CAMLine_132_io_we),
    .io_wi(CAMLine_132_io_wi),
    .io_key(CAMLine_132_io_key),
    .io_din(CAMLine_132_io_din),
    .io_hit(CAMLine_132_io_hit)
  );
  CAMLine CAMLine_133 ( // @[cam.scala 81:36]
    .clock(CAMLine_133_clock),
    .io_we(CAMLine_133_io_we),
    .io_wi(CAMLine_133_io_wi),
    .io_key(CAMLine_133_io_key),
    .io_din(CAMLine_133_io_din),
    .io_hit(CAMLine_133_io_hit)
  );
  CAMLine CAMLine_134 ( // @[cam.scala 81:36]
    .clock(CAMLine_134_clock),
    .io_we(CAMLine_134_io_we),
    .io_wi(CAMLine_134_io_wi),
    .io_key(CAMLine_134_io_key),
    .io_din(CAMLine_134_io_din),
    .io_hit(CAMLine_134_io_hit)
  );
  CAMLine CAMLine_135 ( // @[cam.scala 81:36]
    .clock(CAMLine_135_clock),
    .io_we(CAMLine_135_io_we),
    .io_wi(CAMLine_135_io_wi),
    .io_key(CAMLine_135_io_key),
    .io_din(CAMLine_135_io_din),
    .io_hit(CAMLine_135_io_hit)
  );
  CAMLine CAMLine_136 ( // @[cam.scala 81:36]
    .clock(CAMLine_136_clock),
    .io_we(CAMLine_136_io_we),
    .io_wi(CAMLine_136_io_wi),
    .io_key(CAMLine_136_io_key),
    .io_din(CAMLine_136_io_din),
    .io_hit(CAMLine_136_io_hit)
  );
  CAMLine CAMLine_137 ( // @[cam.scala 81:36]
    .clock(CAMLine_137_clock),
    .io_we(CAMLine_137_io_we),
    .io_wi(CAMLine_137_io_wi),
    .io_key(CAMLine_137_io_key),
    .io_din(CAMLine_137_io_din),
    .io_hit(CAMLine_137_io_hit)
  );
  CAMLine CAMLine_138 ( // @[cam.scala 81:36]
    .clock(CAMLine_138_clock),
    .io_we(CAMLine_138_io_we),
    .io_wi(CAMLine_138_io_wi),
    .io_key(CAMLine_138_io_key),
    .io_din(CAMLine_138_io_din),
    .io_hit(CAMLine_138_io_hit)
  );
  CAMLine CAMLine_139 ( // @[cam.scala 81:36]
    .clock(CAMLine_139_clock),
    .io_we(CAMLine_139_io_we),
    .io_wi(CAMLine_139_io_wi),
    .io_key(CAMLine_139_io_key),
    .io_din(CAMLine_139_io_din),
    .io_hit(CAMLine_139_io_hit)
  );
  CAMLine CAMLine_140 ( // @[cam.scala 81:36]
    .clock(CAMLine_140_clock),
    .io_we(CAMLine_140_io_we),
    .io_wi(CAMLine_140_io_wi),
    .io_key(CAMLine_140_io_key),
    .io_din(CAMLine_140_io_din),
    .io_hit(CAMLine_140_io_hit)
  );
  CAMLine CAMLine_141 ( // @[cam.scala 81:36]
    .clock(CAMLine_141_clock),
    .io_we(CAMLine_141_io_we),
    .io_wi(CAMLine_141_io_wi),
    .io_key(CAMLine_141_io_key),
    .io_din(CAMLine_141_io_din),
    .io_hit(CAMLine_141_io_hit)
  );
  CAMLine CAMLine_142 ( // @[cam.scala 81:36]
    .clock(CAMLine_142_clock),
    .io_we(CAMLine_142_io_we),
    .io_wi(CAMLine_142_io_wi),
    .io_key(CAMLine_142_io_key),
    .io_din(CAMLine_142_io_din),
    .io_hit(CAMLine_142_io_hit)
  );
  CAMLine CAMLine_143 ( // @[cam.scala 81:36]
    .clock(CAMLine_143_clock),
    .io_we(CAMLine_143_io_we),
    .io_wi(CAMLine_143_io_wi),
    .io_key(CAMLine_143_io_key),
    .io_din(CAMLine_143_io_din),
    .io_hit(CAMLine_143_io_hit)
  );
  CAMLine CAMLine_144 ( // @[cam.scala 81:36]
    .clock(CAMLine_144_clock),
    .io_we(CAMLine_144_io_we),
    .io_wi(CAMLine_144_io_wi),
    .io_key(CAMLine_144_io_key),
    .io_din(CAMLine_144_io_din),
    .io_hit(CAMLine_144_io_hit)
  );
  CAMLine CAMLine_145 ( // @[cam.scala 81:36]
    .clock(CAMLine_145_clock),
    .io_we(CAMLine_145_io_we),
    .io_wi(CAMLine_145_io_wi),
    .io_key(CAMLine_145_io_key),
    .io_din(CAMLine_145_io_din),
    .io_hit(CAMLine_145_io_hit)
  );
  CAMLine CAMLine_146 ( // @[cam.scala 81:36]
    .clock(CAMLine_146_clock),
    .io_we(CAMLine_146_io_we),
    .io_wi(CAMLine_146_io_wi),
    .io_key(CAMLine_146_io_key),
    .io_din(CAMLine_146_io_din),
    .io_hit(CAMLine_146_io_hit)
  );
  CAMLine CAMLine_147 ( // @[cam.scala 81:36]
    .clock(CAMLine_147_clock),
    .io_we(CAMLine_147_io_we),
    .io_wi(CAMLine_147_io_wi),
    .io_key(CAMLine_147_io_key),
    .io_din(CAMLine_147_io_din),
    .io_hit(CAMLine_147_io_hit)
  );
  CAMLine CAMLine_148 ( // @[cam.scala 81:36]
    .clock(CAMLine_148_clock),
    .io_we(CAMLine_148_io_we),
    .io_wi(CAMLine_148_io_wi),
    .io_key(CAMLine_148_io_key),
    .io_din(CAMLine_148_io_din),
    .io_hit(CAMLine_148_io_hit)
  );
  CAMLine CAMLine_149 ( // @[cam.scala 81:36]
    .clock(CAMLine_149_clock),
    .io_we(CAMLine_149_io_we),
    .io_wi(CAMLine_149_io_wi),
    .io_key(CAMLine_149_io_key),
    .io_din(CAMLine_149_io_din),
    .io_hit(CAMLine_149_io_hit)
  );
  CAMLine CAMLine_150 ( // @[cam.scala 81:36]
    .clock(CAMLine_150_clock),
    .io_we(CAMLine_150_io_we),
    .io_wi(CAMLine_150_io_wi),
    .io_key(CAMLine_150_io_key),
    .io_din(CAMLine_150_io_din),
    .io_hit(CAMLine_150_io_hit)
  );
  CAMLine CAMLine_151 ( // @[cam.scala 81:36]
    .clock(CAMLine_151_clock),
    .io_we(CAMLine_151_io_we),
    .io_wi(CAMLine_151_io_wi),
    .io_key(CAMLine_151_io_key),
    .io_din(CAMLine_151_io_din),
    .io_hit(CAMLine_151_io_hit)
  );
  CAMLine CAMLine_152 ( // @[cam.scala 81:36]
    .clock(CAMLine_152_clock),
    .io_we(CAMLine_152_io_we),
    .io_wi(CAMLine_152_io_wi),
    .io_key(CAMLine_152_io_key),
    .io_din(CAMLine_152_io_din),
    .io_hit(CAMLine_152_io_hit)
  );
  CAMLine CAMLine_153 ( // @[cam.scala 81:36]
    .clock(CAMLine_153_clock),
    .io_we(CAMLine_153_io_we),
    .io_wi(CAMLine_153_io_wi),
    .io_key(CAMLine_153_io_key),
    .io_din(CAMLine_153_io_din),
    .io_hit(CAMLine_153_io_hit)
  );
  CAMLine CAMLine_154 ( // @[cam.scala 81:36]
    .clock(CAMLine_154_clock),
    .io_we(CAMLine_154_io_we),
    .io_wi(CAMLine_154_io_wi),
    .io_key(CAMLine_154_io_key),
    .io_din(CAMLine_154_io_din),
    .io_hit(CAMLine_154_io_hit)
  );
  CAMLine CAMLine_155 ( // @[cam.scala 81:36]
    .clock(CAMLine_155_clock),
    .io_we(CAMLine_155_io_we),
    .io_wi(CAMLine_155_io_wi),
    .io_key(CAMLine_155_io_key),
    .io_din(CAMLine_155_io_din),
    .io_hit(CAMLine_155_io_hit)
  );
  CAMLine CAMLine_156 ( // @[cam.scala 81:36]
    .clock(CAMLine_156_clock),
    .io_we(CAMLine_156_io_we),
    .io_wi(CAMLine_156_io_wi),
    .io_key(CAMLine_156_io_key),
    .io_din(CAMLine_156_io_din),
    .io_hit(CAMLine_156_io_hit)
  );
  CAMLine CAMLine_157 ( // @[cam.scala 81:36]
    .clock(CAMLine_157_clock),
    .io_we(CAMLine_157_io_we),
    .io_wi(CAMLine_157_io_wi),
    .io_key(CAMLine_157_io_key),
    .io_din(CAMLine_157_io_din),
    .io_hit(CAMLine_157_io_hit)
  );
  CAMLine CAMLine_158 ( // @[cam.scala 81:36]
    .clock(CAMLine_158_clock),
    .io_we(CAMLine_158_io_we),
    .io_wi(CAMLine_158_io_wi),
    .io_key(CAMLine_158_io_key),
    .io_din(CAMLine_158_io_din),
    .io_hit(CAMLine_158_io_hit)
  );
  CAMLine CAMLine_159 ( // @[cam.scala 81:36]
    .clock(CAMLine_159_clock),
    .io_we(CAMLine_159_io_we),
    .io_wi(CAMLine_159_io_wi),
    .io_key(CAMLine_159_io_key),
    .io_din(CAMLine_159_io_din),
    .io_hit(CAMLine_159_io_hit)
  );
  CAMLine CAMLine_160 ( // @[cam.scala 81:36]
    .clock(CAMLine_160_clock),
    .io_we(CAMLine_160_io_we),
    .io_wi(CAMLine_160_io_wi),
    .io_key(CAMLine_160_io_key),
    .io_din(CAMLine_160_io_din),
    .io_hit(CAMLine_160_io_hit)
  );
  CAMLine CAMLine_161 ( // @[cam.scala 81:36]
    .clock(CAMLine_161_clock),
    .io_we(CAMLine_161_io_we),
    .io_wi(CAMLine_161_io_wi),
    .io_key(CAMLine_161_io_key),
    .io_din(CAMLine_161_io_din),
    .io_hit(CAMLine_161_io_hit)
  );
  CAMLine CAMLine_162 ( // @[cam.scala 81:36]
    .clock(CAMLine_162_clock),
    .io_we(CAMLine_162_io_we),
    .io_wi(CAMLine_162_io_wi),
    .io_key(CAMLine_162_io_key),
    .io_din(CAMLine_162_io_din),
    .io_hit(CAMLine_162_io_hit)
  );
  CAMLine CAMLine_163 ( // @[cam.scala 81:36]
    .clock(CAMLine_163_clock),
    .io_we(CAMLine_163_io_we),
    .io_wi(CAMLine_163_io_wi),
    .io_key(CAMLine_163_io_key),
    .io_din(CAMLine_163_io_din),
    .io_hit(CAMLine_163_io_hit)
  );
  CAMLine CAMLine_164 ( // @[cam.scala 81:36]
    .clock(CAMLine_164_clock),
    .io_we(CAMLine_164_io_we),
    .io_wi(CAMLine_164_io_wi),
    .io_key(CAMLine_164_io_key),
    .io_din(CAMLine_164_io_din),
    .io_hit(CAMLine_164_io_hit)
  );
  CAMLine CAMLine_165 ( // @[cam.scala 81:36]
    .clock(CAMLine_165_clock),
    .io_we(CAMLine_165_io_we),
    .io_wi(CAMLine_165_io_wi),
    .io_key(CAMLine_165_io_key),
    .io_din(CAMLine_165_io_din),
    .io_hit(CAMLine_165_io_hit)
  );
  CAMLine CAMLine_166 ( // @[cam.scala 81:36]
    .clock(CAMLine_166_clock),
    .io_we(CAMLine_166_io_we),
    .io_wi(CAMLine_166_io_wi),
    .io_key(CAMLine_166_io_key),
    .io_din(CAMLine_166_io_din),
    .io_hit(CAMLine_166_io_hit)
  );
  CAMLine CAMLine_167 ( // @[cam.scala 81:36]
    .clock(CAMLine_167_clock),
    .io_we(CAMLine_167_io_we),
    .io_wi(CAMLine_167_io_wi),
    .io_key(CAMLine_167_io_key),
    .io_din(CAMLine_167_io_din),
    .io_hit(CAMLine_167_io_hit)
  );
  CAMLine CAMLine_168 ( // @[cam.scala 81:36]
    .clock(CAMLine_168_clock),
    .io_we(CAMLine_168_io_we),
    .io_wi(CAMLine_168_io_wi),
    .io_key(CAMLine_168_io_key),
    .io_din(CAMLine_168_io_din),
    .io_hit(CAMLine_168_io_hit)
  );
  CAMLine CAMLine_169 ( // @[cam.scala 81:36]
    .clock(CAMLine_169_clock),
    .io_we(CAMLine_169_io_we),
    .io_wi(CAMLine_169_io_wi),
    .io_key(CAMLine_169_io_key),
    .io_din(CAMLine_169_io_din),
    .io_hit(CAMLine_169_io_hit)
  );
  CAMLine CAMLine_170 ( // @[cam.scala 81:36]
    .clock(CAMLine_170_clock),
    .io_we(CAMLine_170_io_we),
    .io_wi(CAMLine_170_io_wi),
    .io_key(CAMLine_170_io_key),
    .io_din(CAMLine_170_io_din),
    .io_hit(CAMLine_170_io_hit)
  );
  CAMLine CAMLine_171 ( // @[cam.scala 81:36]
    .clock(CAMLine_171_clock),
    .io_we(CAMLine_171_io_we),
    .io_wi(CAMLine_171_io_wi),
    .io_key(CAMLine_171_io_key),
    .io_din(CAMLine_171_io_din),
    .io_hit(CAMLine_171_io_hit)
  );
  CAMLine CAMLine_172 ( // @[cam.scala 81:36]
    .clock(CAMLine_172_clock),
    .io_we(CAMLine_172_io_we),
    .io_wi(CAMLine_172_io_wi),
    .io_key(CAMLine_172_io_key),
    .io_din(CAMLine_172_io_din),
    .io_hit(CAMLine_172_io_hit)
  );
  CAMLine CAMLine_173 ( // @[cam.scala 81:36]
    .clock(CAMLine_173_clock),
    .io_we(CAMLine_173_io_we),
    .io_wi(CAMLine_173_io_wi),
    .io_key(CAMLine_173_io_key),
    .io_din(CAMLine_173_io_din),
    .io_hit(CAMLine_173_io_hit)
  );
  CAMLine CAMLine_174 ( // @[cam.scala 81:36]
    .clock(CAMLine_174_clock),
    .io_we(CAMLine_174_io_we),
    .io_wi(CAMLine_174_io_wi),
    .io_key(CAMLine_174_io_key),
    .io_din(CAMLine_174_io_din),
    .io_hit(CAMLine_174_io_hit)
  );
  CAMLine CAMLine_175 ( // @[cam.scala 81:36]
    .clock(CAMLine_175_clock),
    .io_we(CAMLine_175_io_we),
    .io_wi(CAMLine_175_io_wi),
    .io_key(CAMLine_175_io_key),
    .io_din(CAMLine_175_io_din),
    .io_hit(CAMLine_175_io_hit)
  );
  CAMLine CAMLine_176 ( // @[cam.scala 81:36]
    .clock(CAMLine_176_clock),
    .io_we(CAMLine_176_io_we),
    .io_wi(CAMLine_176_io_wi),
    .io_key(CAMLine_176_io_key),
    .io_din(CAMLine_176_io_din),
    .io_hit(CAMLine_176_io_hit)
  );
  CAMLine CAMLine_177 ( // @[cam.scala 81:36]
    .clock(CAMLine_177_clock),
    .io_we(CAMLine_177_io_we),
    .io_wi(CAMLine_177_io_wi),
    .io_key(CAMLine_177_io_key),
    .io_din(CAMLine_177_io_din),
    .io_hit(CAMLine_177_io_hit)
  );
  CAMLine CAMLine_178 ( // @[cam.scala 81:36]
    .clock(CAMLine_178_clock),
    .io_we(CAMLine_178_io_we),
    .io_wi(CAMLine_178_io_wi),
    .io_key(CAMLine_178_io_key),
    .io_din(CAMLine_178_io_din),
    .io_hit(CAMLine_178_io_hit)
  );
  CAMLine CAMLine_179 ( // @[cam.scala 81:36]
    .clock(CAMLine_179_clock),
    .io_we(CAMLine_179_io_we),
    .io_wi(CAMLine_179_io_wi),
    .io_key(CAMLine_179_io_key),
    .io_din(CAMLine_179_io_din),
    .io_hit(CAMLine_179_io_hit)
  );
  CAMLine CAMLine_180 ( // @[cam.scala 81:36]
    .clock(CAMLine_180_clock),
    .io_we(CAMLine_180_io_we),
    .io_wi(CAMLine_180_io_wi),
    .io_key(CAMLine_180_io_key),
    .io_din(CAMLine_180_io_din),
    .io_hit(CAMLine_180_io_hit)
  );
  CAMLine CAMLine_181 ( // @[cam.scala 81:36]
    .clock(CAMLine_181_clock),
    .io_we(CAMLine_181_io_we),
    .io_wi(CAMLine_181_io_wi),
    .io_key(CAMLine_181_io_key),
    .io_din(CAMLine_181_io_din),
    .io_hit(CAMLine_181_io_hit)
  );
  CAMLine CAMLine_182 ( // @[cam.scala 81:36]
    .clock(CAMLine_182_clock),
    .io_we(CAMLine_182_io_we),
    .io_wi(CAMLine_182_io_wi),
    .io_key(CAMLine_182_io_key),
    .io_din(CAMLine_182_io_din),
    .io_hit(CAMLine_182_io_hit)
  );
  CAMLine CAMLine_183 ( // @[cam.scala 81:36]
    .clock(CAMLine_183_clock),
    .io_we(CAMLine_183_io_we),
    .io_wi(CAMLine_183_io_wi),
    .io_key(CAMLine_183_io_key),
    .io_din(CAMLine_183_io_din),
    .io_hit(CAMLine_183_io_hit)
  );
  CAMLine CAMLine_184 ( // @[cam.scala 81:36]
    .clock(CAMLine_184_clock),
    .io_we(CAMLine_184_io_we),
    .io_wi(CAMLine_184_io_wi),
    .io_key(CAMLine_184_io_key),
    .io_din(CAMLine_184_io_din),
    .io_hit(CAMLine_184_io_hit)
  );
  CAMLine CAMLine_185 ( // @[cam.scala 81:36]
    .clock(CAMLine_185_clock),
    .io_we(CAMLine_185_io_we),
    .io_wi(CAMLine_185_io_wi),
    .io_key(CAMLine_185_io_key),
    .io_din(CAMLine_185_io_din),
    .io_hit(CAMLine_185_io_hit)
  );
  CAMLine CAMLine_186 ( // @[cam.scala 81:36]
    .clock(CAMLine_186_clock),
    .io_we(CAMLine_186_io_we),
    .io_wi(CAMLine_186_io_wi),
    .io_key(CAMLine_186_io_key),
    .io_din(CAMLine_186_io_din),
    .io_hit(CAMLine_186_io_hit)
  );
  CAMLine CAMLine_187 ( // @[cam.scala 81:36]
    .clock(CAMLine_187_clock),
    .io_we(CAMLine_187_io_we),
    .io_wi(CAMLine_187_io_wi),
    .io_key(CAMLine_187_io_key),
    .io_din(CAMLine_187_io_din),
    .io_hit(CAMLine_187_io_hit)
  );
  CAMLine CAMLine_188 ( // @[cam.scala 81:36]
    .clock(CAMLine_188_clock),
    .io_we(CAMLine_188_io_we),
    .io_wi(CAMLine_188_io_wi),
    .io_key(CAMLine_188_io_key),
    .io_din(CAMLine_188_io_din),
    .io_hit(CAMLine_188_io_hit)
  );
  CAMLine CAMLine_189 ( // @[cam.scala 81:36]
    .clock(CAMLine_189_clock),
    .io_we(CAMLine_189_io_we),
    .io_wi(CAMLine_189_io_wi),
    .io_key(CAMLine_189_io_key),
    .io_din(CAMLine_189_io_din),
    .io_hit(CAMLine_189_io_hit)
  );
  CAMLine CAMLine_190 ( // @[cam.scala 81:36]
    .clock(CAMLine_190_clock),
    .io_we(CAMLine_190_io_we),
    .io_wi(CAMLine_190_io_wi),
    .io_key(CAMLine_190_io_key),
    .io_din(CAMLine_190_io_din),
    .io_hit(CAMLine_190_io_hit)
  );
  CAMLine CAMLine_191 ( // @[cam.scala 81:36]
    .clock(CAMLine_191_clock),
    .io_we(CAMLine_191_io_we),
    .io_wi(CAMLine_191_io_wi),
    .io_key(CAMLine_191_io_key),
    .io_din(CAMLine_191_io_din),
    .io_hit(CAMLine_191_io_hit)
  );
  CAMLine CAMLine_192 ( // @[cam.scala 81:36]
    .clock(CAMLine_192_clock),
    .io_we(CAMLine_192_io_we),
    .io_wi(CAMLine_192_io_wi),
    .io_key(CAMLine_192_io_key),
    .io_din(CAMLine_192_io_din),
    .io_hit(CAMLine_192_io_hit)
  );
  CAMLine CAMLine_193 ( // @[cam.scala 81:36]
    .clock(CAMLine_193_clock),
    .io_we(CAMLine_193_io_we),
    .io_wi(CAMLine_193_io_wi),
    .io_key(CAMLine_193_io_key),
    .io_din(CAMLine_193_io_din),
    .io_hit(CAMLine_193_io_hit)
  );
  CAMLine CAMLine_194 ( // @[cam.scala 81:36]
    .clock(CAMLine_194_clock),
    .io_we(CAMLine_194_io_we),
    .io_wi(CAMLine_194_io_wi),
    .io_key(CAMLine_194_io_key),
    .io_din(CAMLine_194_io_din),
    .io_hit(CAMLine_194_io_hit)
  );
  CAMLine CAMLine_195 ( // @[cam.scala 81:36]
    .clock(CAMLine_195_clock),
    .io_we(CAMLine_195_io_we),
    .io_wi(CAMLine_195_io_wi),
    .io_key(CAMLine_195_io_key),
    .io_din(CAMLine_195_io_din),
    .io_hit(CAMLine_195_io_hit)
  );
  CAMLine CAMLine_196 ( // @[cam.scala 81:36]
    .clock(CAMLine_196_clock),
    .io_we(CAMLine_196_io_we),
    .io_wi(CAMLine_196_io_wi),
    .io_key(CAMLine_196_io_key),
    .io_din(CAMLine_196_io_din),
    .io_hit(CAMLine_196_io_hit)
  );
  CAMLine CAMLine_197 ( // @[cam.scala 81:36]
    .clock(CAMLine_197_clock),
    .io_we(CAMLine_197_io_we),
    .io_wi(CAMLine_197_io_wi),
    .io_key(CAMLine_197_io_key),
    .io_din(CAMLine_197_io_din),
    .io_hit(CAMLine_197_io_hit)
  );
  CAMLine CAMLine_198 ( // @[cam.scala 81:36]
    .clock(CAMLine_198_clock),
    .io_we(CAMLine_198_io_we),
    .io_wi(CAMLine_198_io_wi),
    .io_key(CAMLine_198_io_key),
    .io_din(CAMLine_198_io_din),
    .io_hit(CAMLine_198_io_hit)
  );
  CAMLine CAMLine_199 ( // @[cam.scala 81:36]
    .clock(CAMLine_199_clock),
    .io_we(CAMLine_199_io_we),
    .io_wi(CAMLine_199_io_wi),
    .io_key(CAMLine_199_io_key),
    .io_din(CAMLine_199_io_din),
    .io_hit(CAMLine_199_io_hit)
  );
  CAMLine CAMLine_200 ( // @[cam.scala 81:36]
    .clock(CAMLine_200_clock),
    .io_we(CAMLine_200_io_we),
    .io_wi(CAMLine_200_io_wi),
    .io_key(CAMLine_200_io_key),
    .io_din(CAMLine_200_io_din),
    .io_hit(CAMLine_200_io_hit)
  );
  CAMLine CAMLine_201 ( // @[cam.scala 81:36]
    .clock(CAMLine_201_clock),
    .io_we(CAMLine_201_io_we),
    .io_wi(CAMLine_201_io_wi),
    .io_key(CAMLine_201_io_key),
    .io_din(CAMLine_201_io_din),
    .io_hit(CAMLine_201_io_hit)
  );
  CAMLine CAMLine_202 ( // @[cam.scala 81:36]
    .clock(CAMLine_202_clock),
    .io_we(CAMLine_202_io_we),
    .io_wi(CAMLine_202_io_wi),
    .io_key(CAMLine_202_io_key),
    .io_din(CAMLine_202_io_din),
    .io_hit(CAMLine_202_io_hit)
  );
  CAMLine CAMLine_203 ( // @[cam.scala 81:36]
    .clock(CAMLine_203_clock),
    .io_we(CAMLine_203_io_we),
    .io_wi(CAMLine_203_io_wi),
    .io_key(CAMLine_203_io_key),
    .io_din(CAMLine_203_io_din),
    .io_hit(CAMLine_203_io_hit)
  );
  CAMLine CAMLine_204 ( // @[cam.scala 81:36]
    .clock(CAMLine_204_clock),
    .io_we(CAMLine_204_io_we),
    .io_wi(CAMLine_204_io_wi),
    .io_key(CAMLine_204_io_key),
    .io_din(CAMLine_204_io_din),
    .io_hit(CAMLine_204_io_hit)
  );
  CAMLine CAMLine_205 ( // @[cam.scala 81:36]
    .clock(CAMLine_205_clock),
    .io_we(CAMLine_205_io_we),
    .io_wi(CAMLine_205_io_wi),
    .io_key(CAMLine_205_io_key),
    .io_din(CAMLine_205_io_din),
    .io_hit(CAMLine_205_io_hit)
  );
  CAMLine CAMLine_206 ( // @[cam.scala 81:36]
    .clock(CAMLine_206_clock),
    .io_we(CAMLine_206_io_we),
    .io_wi(CAMLine_206_io_wi),
    .io_key(CAMLine_206_io_key),
    .io_din(CAMLine_206_io_din),
    .io_hit(CAMLine_206_io_hit)
  );
  CAMLine CAMLine_207 ( // @[cam.scala 81:36]
    .clock(CAMLine_207_clock),
    .io_we(CAMLine_207_io_we),
    .io_wi(CAMLine_207_io_wi),
    .io_key(CAMLine_207_io_key),
    .io_din(CAMLine_207_io_din),
    .io_hit(CAMLine_207_io_hit)
  );
  CAMLine CAMLine_208 ( // @[cam.scala 81:36]
    .clock(CAMLine_208_clock),
    .io_we(CAMLine_208_io_we),
    .io_wi(CAMLine_208_io_wi),
    .io_key(CAMLine_208_io_key),
    .io_din(CAMLine_208_io_din),
    .io_hit(CAMLine_208_io_hit)
  );
  CAMLine CAMLine_209 ( // @[cam.scala 81:36]
    .clock(CAMLine_209_clock),
    .io_we(CAMLine_209_io_we),
    .io_wi(CAMLine_209_io_wi),
    .io_key(CAMLine_209_io_key),
    .io_din(CAMLine_209_io_din),
    .io_hit(CAMLine_209_io_hit)
  );
  CAMLine CAMLine_210 ( // @[cam.scala 81:36]
    .clock(CAMLine_210_clock),
    .io_we(CAMLine_210_io_we),
    .io_wi(CAMLine_210_io_wi),
    .io_key(CAMLine_210_io_key),
    .io_din(CAMLine_210_io_din),
    .io_hit(CAMLine_210_io_hit)
  );
  CAMLine CAMLine_211 ( // @[cam.scala 81:36]
    .clock(CAMLine_211_clock),
    .io_we(CAMLine_211_io_we),
    .io_wi(CAMLine_211_io_wi),
    .io_key(CAMLine_211_io_key),
    .io_din(CAMLine_211_io_din),
    .io_hit(CAMLine_211_io_hit)
  );
  CAMLine CAMLine_212 ( // @[cam.scala 81:36]
    .clock(CAMLine_212_clock),
    .io_we(CAMLine_212_io_we),
    .io_wi(CAMLine_212_io_wi),
    .io_key(CAMLine_212_io_key),
    .io_din(CAMLine_212_io_din),
    .io_hit(CAMLine_212_io_hit)
  );
  CAMLine CAMLine_213 ( // @[cam.scala 81:36]
    .clock(CAMLine_213_clock),
    .io_we(CAMLine_213_io_we),
    .io_wi(CAMLine_213_io_wi),
    .io_key(CAMLine_213_io_key),
    .io_din(CAMLine_213_io_din),
    .io_hit(CAMLine_213_io_hit)
  );
  CAMLine CAMLine_214 ( // @[cam.scala 81:36]
    .clock(CAMLine_214_clock),
    .io_we(CAMLine_214_io_we),
    .io_wi(CAMLine_214_io_wi),
    .io_key(CAMLine_214_io_key),
    .io_din(CAMLine_214_io_din),
    .io_hit(CAMLine_214_io_hit)
  );
  CAMLine CAMLine_215 ( // @[cam.scala 81:36]
    .clock(CAMLine_215_clock),
    .io_we(CAMLine_215_io_we),
    .io_wi(CAMLine_215_io_wi),
    .io_key(CAMLine_215_io_key),
    .io_din(CAMLine_215_io_din),
    .io_hit(CAMLine_215_io_hit)
  );
  CAMLine CAMLine_216 ( // @[cam.scala 81:36]
    .clock(CAMLine_216_clock),
    .io_we(CAMLine_216_io_we),
    .io_wi(CAMLine_216_io_wi),
    .io_key(CAMLine_216_io_key),
    .io_din(CAMLine_216_io_din),
    .io_hit(CAMLine_216_io_hit)
  );
  CAMLine CAMLine_217 ( // @[cam.scala 81:36]
    .clock(CAMLine_217_clock),
    .io_we(CAMLine_217_io_we),
    .io_wi(CAMLine_217_io_wi),
    .io_key(CAMLine_217_io_key),
    .io_din(CAMLine_217_io_din),
    .io_hit(CAMLine_217_io_hit)
  );
  CAMLine CAMLine_218 ( // @[cam.scala 81:36]
    .clock(CAMLine_218_clock),
    .io_we(CAMLine_218_io_we),
    .io_wi(CAMLine_218_io_wi),
    .io_key(CAMLine_218_io_key),
    .io_din(CAMLine_218_io_din),
    .io_hit(CAMLine_218_io_hit)
  );
  CAMLine CAMLine_219 ( // @[cam.scala 81:36]
    .clock(CAMLine_219_clock),
    .io_we(CAMLine_219_io_we),
    .io_wi(CAMLine_219_io_wi),
    .io_key(CAMLine_219_io_key),
    .io_din(CAMLine_219_io_din),
    .io_hit(CAMLine_219_io_hit)
  );
  CAMLine CAMLine_220 ( // @[cam.scala 81:36]
    .clock(CAMLine_220_clock),
    .io_we(CAMLine_220_io_we),
    .io_wi(CAMLine_220_io_wi),
    .io_key(CAMLine_220_io_key),
    .io_din(CAMLine_220_io_din),
    .io_hit(CAMLine_220_io_hit)
  );
  CAMLine CAMLine_221 ( // @[cam.scala 81:36]
    .clock(CAMLine_221_clock),
    .io_we(CAMLine_221_io_we),
    .io_wi(CAMLine_221_io_wi),
    .io_key(CAMLine_221_io_key),
    .io_din(CAMLine_221_io_din),
    .io_hit(CAMLine_221_io_hit)
  );
  CAMLine CAMLine_222 ( // @[cam.scala 81:36]
    .clock(CAMLine_222_clock),
    .io_we(CAMLine_222_io_we),
    .io_wi(CAMLine_222_io_wi),
    .io_key(CAMLine_222_io_key),
    .io_din(CAMLine_222_io_din),
    .io_hit(CAMLine_222_io_hit)
  );
  CAMLine CAMLine_223 ( // @[cam.scala 81:36]
    .clock(CAMLine_223_clock),
    .io_we(CAMLine_223_io_we),
    .io_wi(CAMLine_223_io_wi),
    .io_key(CAMLine_223_io_key),
    .io_din(CAMLine_223_io_din),
    .io_hit(CAMLine_223_io_hit)
  );
  CAMLine CAMLine_224 ( // @[cam.scala 81:36]
    .clock(CAMLine_224_clock),
    .io_we(CAMLine_224_io_we),
    .io_wi(CAMLine_224_io_wi),
    .io_key(CAMLine_224_io_key),
    .io_din(CAMLine_224_io_din),
    .io_hit(CAMLine_224_io_hit)
  );
  CAMLine CAMLine_225 ( // @[cam.scala 81:36]
    .clock(CAMLine_225_clock),
    .io_we(CAMLine_225_io_we),
    .io_wi(CAMLine_225_io_wi),
    .io_key(CAMLine_225_io_key),
    .io_din(CAMLine_225_io_din),
    .io_hit(CAMLine_225_io_hit)
  );
  CAMLine CAMLine_226 ( // @[cam.scala 81:36]
    .clock(CAMLine_226_clock),
    .io_we(CAMLine_226_io_we),
    .io_wi(CAMLine_226_io_wi),
    .io_key(CAMLine_226_io_key),
    .io_din(CAMLine_226_io_din),
    .io_hit(CAMLine_226_io_hit)
  );
  CAMLine CAMLine_227 ( // @[cam.scala 81:36]
    .clock(CAMLine_227_clock),
    .io_we(CAMLine_227_io_we),
    .io_wi(CAMLine_227_io_wi),
    .io_key(CAMLine_227_io_key),
    .io_din(CAMLine_227_io_din),
    .io_hit(CAMLine_227_io_hit)
  );
  CAMLine CAMLine_228 ( // @[cam.scala 81:36]
    .clock(CAMLine_228_clock),
    .io_we(CAMLine_228_io_we),
    .io_wi(CAMLine_228_io_wi),
    .io_key(CAMLine_228_io_key),
    .io_din(CAMLine_228_io_din),
    .io_hit(CAMLine_228_io_hit)
  );
  CAMLine CAMLine_229 ( // @[cam.scala 81:36]
    .clock(CAMLine_229_clock),
    .io_we(CAMLine_229_io_we),
    .io_wi(CAMLine_229_io_wi),
    .io_key(CAMLine_229_io_key),
    .io_din(CAMLine_229_io_din),
    .io_hit(CAMLine_229_io_hit)
  );
  CAMLine CAMLine_230 ( // @[cam.scala 81:36]
    .clock(CAMLine_230_clock),
    .io_we(CAMLine_230_io_we),
    .io_wi(CAMLine_230_io_wi),
    .io_key(CAMLine_230_io_key),
    .io_din(CAMLine_230_io_din),
    .io_hit(CAMLine_230_io_hit)
  );
  CAMLine CAMLine_231 ( // @[cam.scala 81:36]
    .clock(CAMLine_231_clock),
    .io_we(CAMLine_231_io_we),
    .io_wi(CAMLine_231_io_wi),
    .io_key(CAMLine_231_io_key),
    .io_din(CAMLine_231_io_din),
    .io_hit(CAMLine_231_io_hit)
  );
  CAMLine CAMLine_232 ( // @[cam.scala 81:36]
    .clock(CAMLine_232_clock),
    .io_we(CAMLine_232_io_we),
    .io_wi(CAMLine_232_io_wi),
    .io_key(CAMLine_232_io_key),
    .io_din(CAMLine_232_io_din),
    .io_hit(CAMLine_232_io_hit)
  );
  CAMLine CAMLine_233 ( // @[cam.scala 81:36]
    .clock(CAMLine_233_clock),
    .io_we(CAMLine_233_io_we),
    .io_wi(CAMLine_233_io_wi),
    .io_key(CAMLine_233_io_key),
    .io_din(CAMLine_233_io_din),
    .io_hit(CAMLine_233_io_hit)
  );
  CAMLine CAMLine_234 ( // @[cam.scala 81:36]
    .clock(CAMLine_234_clock),
    .io_we(CAMLine_234_io_we),
    .io_wi(CAMLine_234_io_wi),
    .io_key(CAMLine_234_io_key),
    .io_din(CAMLine_234_io_din),
    .io_hit(CAMLine_234_io_hit)
  );
  CAMLine CAMLine_235 ( // @[cam.scala 81:36]
    .clock(CAMLine_235_clock),
    .io_we(CAMLine_235_io_we),
    .io_wi(CAMLine_235_io_wi),
    .io_key(CAMLine_235_io_key),
    .io_din(CAMLine_235_io_din),
    .io_hit(CAMLine_235_io_hit)
  );
  CAMLine CAMLine_236 ( // @[cam.scala 81:36]
    .clock(CAMLine_236_clock),
    .io_we(CAMLine_236_io_we),
    .io_wi(CAMLine_236_io_wi),
    .io_key(CAMLine_236_io_key),
    .io_din(CAMLine_236_io_din),
    .io_hit(CAMLine_236_io_hit)
  );
  CAMLine CAMLine_237 ( // @[cam.scala 81:36]
    .clock(CAMLine_237_clock),
    .io_we(CAMLine_237_io_we),
    .io_wi(CAMLine_237_io_wi),
    .io_key(CAMLine_237_io_key),
    .io_din(CAMLine_237_io_din),
    .io_hit(CAMLine_237_io_hit)
  );
  CAMLine CAMLine_238 ( // @[cam.scala 81:36]
    .clock(CAMLine_238_clock),
    .io_we(CAMLine_238_io_we),
    .io_wi(CAMLine_238_io_wi),
    .io_key(CAMLine_238_io_key),
    .io_din(CAMLine_238_io_din),
    .io_hit(CAMLine_238_io_hit)
  );
  CAMLine CAMLine_239 ( // @[cam.scala 81:36]
    .clock(CAMLine_239_clock),
    .io_we(CAMLine_239_io_we),
    .io_wi(CAMLine_239_io_wi),
    .io_key(CAMLine_239_io_key),
    .io_din(CAMLine_239_io_din),
    .io_hit(CAMLine_239_io_hit)
  );
  CAMLine CAMLine_240 ( // @[cam.scala 81:36]
    .clock(CAMLine_240_clock),
    .io_we(CAMLine_240_io_we),
    .io_wi(CAMLine_240_io_wi),
    .io_key(CAMLine_240_io_key),
    .io_din(CAMLine_240_io_din),
    .io_hit(CAMLine_240_io_hit)
  );
  CAMLine CAMLine_241 ( // @[cam.scala 81:36]
    .clock(CAMLine_241_clock),
    .io_we(CAMLine_241_io_we),
    .io_wi(CAMLine_241_io_wi),
    .io_key(CAMLine_241_io_key),
    .io_din(CAMLine_241_io_din),
    .io_hit(CAMLine_241_io_hit)
  );
  CAMLine CAMLine_242 ( // @[cam.scala 81:36]
    .clock(CAMLine_242_clock),
    .io_we(CAMLine_242_io_we),
    .io_wi(CAMLine_242_io_wi),
    .io_key(CAMLine_242_io_key),
    .io_din(CAMLine_242_io_din),
    .io_hit(CAMLine_242_io_hit)
  );
  CAMLine CAMLine_243 ( // @[cam.scala 81:36]
    .clock(CAMLine_243_clock),
    .io_we(CAMLine_243_io_we),
    .io_wi(CAMLine_243_io_wi),
    .io_key(CAMLine_243_io_key),
    .io_din(CAMLine_243_io_din),
    .io_hit(CAMLine_243_io_hit)
  );
  CAMLine CAMLine_244 ( // @[cam.scala 81:36]
    .clock(CAMLine_244_clock),
    .io_we(CAMLine_244_io_we),
    .io_wi(CAMLine_244_io_wi),
    .io_key(CAMLine_244_io_key),
    .io_din(CAMLine_244_io_din),
    .io_hit(CAMLine_244_io_hit)
  );
  CAMLine CAMLine_245 ( // @[cam.scala 81:36]
    .clock(CAMLine_245_clock),
    .io_we(CAMLine_245_io_we),
    .io_wi(CAMLine_245_io_wi),
    .io_key(CAMLine_245_io_key),
    .io_din(CAMLine_245_io_din),
    .io_hit(CAMLine_245_io_hit)
  );
  CAMLine CAMLine_246 ( // @[cam.scala 81:36]
    .clock(CAMLine_246_clock),
    .io_we(CAMLine_246_io_we),
    .io_wi(CAMLine_246_io_wi),
    .io_key(CAMLine_246_io_key),
    .io_din(CAMLine_246_io_din),
    .io_hit(CAMLine_246_io_hit)
  );
  CAMLine CAMLine_247 ( // @[cam.scala 81:36]
    .clock(CAMLine_247_clock),
    .io_we(CAMLine_247_io_we),
    .io_wi(CAMLine_247_io_wi),
    .io_key(CAMLine_247_io_key),
    .io_din(CAMLine_247_io_din),
    .io_hit(CAMLine_247_io_hit)
  );
  CAMLine CAMLine_248 ( // @[cam.scala 81:36]
    .clock(CAMLine_248_clock),
    .io_we(CAMLine_248_io_we),
    .io_wi(CAMLine_248_io_wi),
    .io_key(CAMLine_248_io_key),
    .io_din(CAMLine_248_io_din),
    .io_hit(CAMLine_248_io_hit)
  );
  CAMLine CAMLine_249 ( // @[cam.scala 81:36]
    .clock(CAMLine_249_clock),
    .io_we(CAMLine_249_io_we),
    .io_wi(CAMLine_249_io_wi),
    .io_key(CAMLine_249_io_key),
    .io_din(CAMLine_249_io_din),
    .io_hit(CAMLine_249_io_hit)
  );
  CAMLine CAMLine_250 ( // @[cam.scala 81:36]
    .clock(CAMLine_250_clock),
    .io_we(CAMLine_250_io_we),
    .io_wi(CAMLine_250_io_wi),
    .io_key(CAMLine_250_io_key),
    .io_din(CAMLine_250_io_din),
    .io_hit(CAMLine_250_io_hit)
  );
  CAMLine CAMLine_251 ( // @[cam.scala 81:36]
    .clock(CAMLine_251_clock),
    .io_we(CAMLine_251_io_we),
    .io_wi(CAMLine_251_io_wi),
    .io_key(CAMLine_251_io_key),
    .io_din(CAMLine_251_io_din),
    .io_hit(CAMLine_251_io_hit)
  );
  CAMLine CAMLine_252 ( // @[cam.scala 81:36]
    .clock(CAMLine_252_clock),
    .io_we(CAMLine_252_io_we),
    .io_wi(CAMLine_252_io_wi),
    .io_key(CAMLine_252_io_key),
    .io_din(CAMLine_252_io_din),
    .io_hit(CAMLine_252_io_hit)
  );
  CAMLine CAMLine_253 ( // @[cam.scala 81:36]
    .clock(CAMLine_253_clock),
    .io_we(CAMLine_253_io_we),
    .io_wi(CAMLine_253_io_wi),
    .io_key(CAMLine_253_io_key),
    .io_din(CAMLine_253_io_din),
    .io_hit(CAMLine_253_io_hit)
  );
  CAMLine CAMLine_254 ( // @[cam.scala 81:36]
    .clock(CAMLine_254_clock),
    .io_we(CAMLine_254_io_we),
    .io_wi(CAMLine_254_io_wi),
    .io_key(CAMLine_254_io_key),
    .io_din(CAMLine_254_io_din),
    .io_hit(CAMLine_254_io_hit)
  );
  CAMLine CAMLine_255 ( // @[cam.scala 81:36]
    .clock(CAMLine_255_clock),
    .io_we(CAMLine_255_io_we),
    .io_wi(CAMLine_255_io_wi),
    .io_key(CAMLine_255_io_key),
    .io_din(CAMLine_255_io_din),
    .io_hit(CAMLine_255_io_hit)
  );
  assign io_hit = _io_hit_T_239 | CAMLine_241_io_hit | CAMLine_242_io_hit | CAMLine_243_io_hit | CAMLine_244_io_hit |
    CAMLine_245_io_hit | CAMLine_246_io_hit | CAMLine_247_io_hit | CAMLine_248_io_hit | CAMLine_249_io_hit |
    CAMLine_250_io_hit | CAMLine_251_io_hit | CAMLine_252_io_hit | CAMLine_253_io_hit | CAMLine_254_io_hit |
    CAMLine_255_io_hit; // @[cam.scala 93:27]
  assign CAMLine_clock = clock;
  assign CAMLine_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_io_wi = io_waddr[0]; // @[cam.scala 86:31]
  assign CAMLine_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_1_clock = clock;
  assign CAMLine_1_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_1_io_wi = io_waddr[1]; // @[cam.scala 86:31]
  assign CAMLine_1_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_1_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_2_clock = clock;
  assign CAMLine_2_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_2_io_wi = io_waddr[2]; // @[cam.scala 86:31]
  assign CAMLine_2_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_2_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_3_clock = clock;
  assign CAMLine_3_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_3_io_wi = io_waddr[3]; // @[cam.scala 86:31]
  assign CAMLine_3_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_3_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_4_clock = clock;
  assign CAMLine_4_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_4_io_wi = io_waddr[4]; // @[cam.scala 86:31]
  assign CAMLine_4_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_4_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_5_clock = clock;
  assign CAMLine_5_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_5_io_wi = io_waddr[5]; // @[cam.scala 86:31]
  assign CAMLine_5_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_5_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_6_clock = clock;
  assign CAMLine_6_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_6_io_wi = io_waddr[6]; // @[cam.scala 86:31]
  assign CAMLine_6_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_6_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_7_clock = clock;
  assign CAMLine_7_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_7_io_wi = io_waddr[7]; // @[cam.scala 86:31]
  assign CAMLine_7_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_7_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_8_clock = clock;
  assign CAMLine_8_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_8_io_wi = io_waddr[8]; // @[cam.scala 86:31]
  assign CAMLine_8_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_8_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_9_clock = clock;
  assign CAMLine_9_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_9_io_wi = io_waddr[9]; // @[cam.scala 86:31]
  assign CAMLine_9_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_9_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_10_clock = clock;
  assign CAMLine_10_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_10_io_wi = io_waddr[10]; // @[cam.scala 86:31]
  assign CAMLine_10_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_10_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_11_clock = clock;
  assign CAMLine_11_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_11_io_wi = io_waddr[11]; // @[cam.scala 86:31]
  assign CAMLine_11_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_11_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_12_clock = clock;
  assign CAMLine_12_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_12_io_wi = io_waddr[12]; // @[cam.scala 86:31]
  assign CAMLine_12_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_12_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_13_clock = clock;
  assign CAMLine_13_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_13_io_wi = io_waddr[13]; // @[cam.scala 86:31]
  assign CAMLine_13_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_13_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_14_clock = clock;
  assign CAMLine_14_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_14_io_wi = io_waddr[14]; // @[cam.scala 86:31]
  assign CAMLine_14_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_14_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_15_clock = clock;
  assign CAMLine_15_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_15_io_wi = io_waddr[15]; // @[cam.scala 86:31]
  assign CAMLine_15_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_15_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_16_clock = clock;
  assign CAMLine_16_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_16_io_wi = io_waddr[16]; // @[cam.scala 86:31]
  assign CAMLine_16_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_16_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_17_clock = clock;
  assign CAMLine_17_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_17_io_wi = io_waddr[17]; // @[cam.scala 86:31]
  assign CAMLine_17_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_17_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_18_clock = clock;
  assign CAMLine_18_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_18_io_wi = io_waddr[18]; // @[cam.scala 86:31]
  assign CAMLine_18_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_18_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_19_clock = clock;
  assign CAMLine_19_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_19_io_wi = io_waddr[19]; // @[cam.scala 86:31]
  assign CAMLine_19_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_19_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_20_clock = clock;
  assign CAMLine_20_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_20_io_wi = io_waddr[20]; // @[cam.scala 86:31]
  assign CAMLine_20_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_20_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_21_clock = clock;
  assign CAMLine_21_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_21_io_wi = io_waddr[21]; // @[cam.scala 86:31]
  assign CAMLine_21_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_21_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_22_clock = clock;
  assign CAMLine_22_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_22_io_wi = io_waddr[22]; // @[cam.scala 86:31]
  assign CAMLine_22_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_22_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_23_clock = clock;
  assign CAMLine_23_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_23_io_wi = io_waddr[23]; // @[cam.scala 86:31]
  assign CAMLine_23_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_23_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_24_clock = clock;
  assign CAMLine_24_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_24_io_wi = io_waddr[24]; // @[cam.scala 86:31]
  assign CAMLine_24_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_24_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_25_clock = clock;
  assign CAMLine_25_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_25_io_wi = io_waddr[25]; // @[cam.scala 86:31]
  assign CAMLine_25_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_25_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_26_clock = clock;
  assign CAMLine_26_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_26_io_wi = io_waddr[26]; // @[cam.scala 86:31]
  assign CAMLine_26_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_26_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_27_clock = clock;
  assign CAMLine_27_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_27_io_wi = io_waddr[27]; // @[cam.scala 86:31]
  assign CAMLine_27_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_27_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_28_clock = clock;
  assign CAMLine_28_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_28_io_wi = io_waddr[28]; // @[cam.scala 86:31]
  assign CAMLine_28_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_28_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_29_clock = clock;
  assign CAMLine_29_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_29_io_wi = io_waddr[29]; // @[cam.scala 86:31]
  assign CAMLine_29_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_29_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_30_clock = clock;
  assign CAMLine_30_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_30_io_wi = io_waddr[30]; // @[cam.scala 86:31]
  assign CAMLine_30_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_30_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_31_clock = clock;
  assign CAMLine_31_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_31_io_wi = io_waddr[31]; // @[cam.scala 86:31]
  assign CAMLine_31_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_31_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_32_clock = clock;
  assign CAMLine_32_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_32_io_wi = io_waddr[32]; // @[cam.scala 86:31]
  assign CAMLine_32_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_32_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_33_clock = clock;
  assign CAMLine_33_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_33_io_wi = io_waddr[33]; // @[cam.scala 86:31]
  assign CAMLine_33_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_33_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_34_clock = clock;
  assign CAMLine_34_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_34_io_wi = io_waddr[34]; // @[cam.scala 86:31]
  assign CAMLine_34_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_34_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_35_clock = clock;
  assign CAMLine_35_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_35_io_wi = io_waddr[35]; // @[cam.scala 86:31]
  assign CAMLine_35_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_35_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_36_clock = clock;
  assign CAMLine_36_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_36_io_wi = io_waddr[36]; // @[cam.scala 86:31]
  assign CAMLine_36_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_36_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_37_clock = clock;
  assign CAMLine_37_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_37_io_wi = io_waddr[37]; // @[cam.scala 86:31]
  assign CAMLine_37_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_37_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_38_clock = clock;
  assign CAMLine_38_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_38_io_wi = io_waddr[38]; // @[cam.scala 86:31]
  assign CAMLine_38_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_38_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_39_clock = clock;
  assign CAMLine_39_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_39_io_wi = io_waddr[39]; // @[cam.scala 86:31]
  assign CAMLine_39_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_39_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_40_clock = clock;
  assign CAMLine_40_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_40_io_wi = io_waddr[40]; // @[cam.scala 86:31]
  assign CAMLine_40_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_40_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_41_clock = clock;
  assign CAMLine_41_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_41_io_wi = io_waddr[41]; // @[cam.scala 86:31]
  assign CAMLine_41_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_41_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_42_clock = clock;
  assign CAMLine_42_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_42_io_wi = io_waddr[42]; // @[cam.scala 86:31]
  assign CAMLine_42_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_42_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_43_clock = clock;
  assign CAMLine_43_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_43_io_wi = io_waddr[43]; // @[cam.scala 86:31]
  assign CAMLine_43_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_43_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_44_clock = clock;
  assign CAMLine_44_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_44_io_wi = io_waddr[44]; // @[cam.scala 86:31]
  assign CAMLine_44_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_44_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_45_clock = clock;
  assign CAMLine_45_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_45_io_wi = io_waddr[45]; // @[cam.scala 86:31]
  assign CAMLine_45_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_45_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_46_clock = clock;
  assign CAMLine_46_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_46_io_wi = io_waddr[46]; // @[cam.scala 86:31]
  assign CAMLine_46_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_46_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_47_clock = clock;
  assign CAMLine_47_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_47_io_wi = io_waddr[47]; // @[cam.scala 86:31]
  assign CAMLine_47_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_47_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_48_clock = clock;
  assign CAMLine_48_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_48_io_wi = io_waddr[48]; // @[cam.scala 86:31]
  assign CAMLine_48_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_48_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_49_clock = clock;
  assign CAMLine_49_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_49_io_wi = io_waddr[49]; // @[cam.scala 86:31]
  assign CAMLine_49_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_49_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_50_clock = clock;
  assign CAMLine_50_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_50_io_wi = io_waddr[50]; // @[cam.scala 86:31]
  assign CAMLine_50_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_50_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_51_clock = clock;
  assign CAMLine_51_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_51_io_wi = io_waddr[51]; // @[cam.scala 86:31]
  assign CAMLine_51_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_51_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_52_clock = clock;
  assign CAMLine_52_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_52_io_wi = io_waddr[52]; // @[cam.scala 86:31]
  assign CAMLine_52_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_52_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_53_clock = clock;
  assign CAMLine_53_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_53_io_wi = io_waddr[53]; // @[cam.scala 86:31]
  assign CAMLine_53_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_53_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_54_clock = clock;
  assign CAMLine_54_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_54_io_wi = io_waddr[54]; // @[cam.scala 86:31]
  assign CAMLine_54_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_54_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_55_clock = clock;
  assign CAMLine_55_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_55_io_wi = io_waddr[55]; // @[cam.scala 86:31]
  assign CAMLine_55_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_55_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_56_clock = clock;
  assign CAMLine_56_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_56_io_wi = io_waddr[56]; // @[cam.scala 86:31]
  assign CAMLine_56_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_56_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_57_clock = clock;
  assign CAMLine_57_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_57_io_wi = io_waddr[57]; // @[cam.scala 86:31]
  assign CAMLine_57_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_57_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_58_clock = clock;
  assign CAMLine_58_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_58_io_wi = io_waddr[58]; // @[cam.scala 86:31]
  assign CAMLine_58_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_58_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_59_clock = clock;
  assign CAMLine_59_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_59_io_wi = io_waddr[59]; // @[cam.scala 86:31]
  assign CAMLine_59_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_59_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_60_clock = clock;
  assign CAMLine_60_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_60_io_wi = io_waddr[60]; // @[cam.scala 86:31]
  assign CAMLine_60_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_60_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_61_clock = clock;
  assign CAMLine_61_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_61_io_wi = io_waddr[61]; // @[cam.scala 86:31]
  assign CAMLine_61_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_61_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_62_clock = clock;
  assign CAMLine_62_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_62_io_wi = io_waddr[62]; // @[cam.scala 86:31]
  assign CAMLine_62_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_62_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_63_clock = clock;
  assign CAMLine_63_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_63_io_wi = io_waddr[63]; // @[cam.scala 86:31]
  assign CAMLine_63_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_63_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_64_clock = clock;
  assign CAMLine_64_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_64_io_wi = io_waddr[64]; // @[cam.scala 86:31]
  assign CAMLine_64_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_64_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_65_clock = clock;
  assign CAMLine_65_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_65_io_wi = io_waddr[65]; // @[cam.scala 86:31]
  assign CAMLine_65_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_65_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_66_clock = clock;
  assign CAMLine_66_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_66_io_wi = io_waddr[66]; // @[cam.scala 86:31]
  assign CAMLine_66_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_66_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_67_clock = clock;
  assign CAMLine_67_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_67_io_wi = io_waddr[67]; // @[cam.scala 86:31]
  assign CAMLine_67_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_67_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_68_clock = clock;
  assign CAMLine_68_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_68_io_wi = io_waddr[68]; // @[cam.scala 86:31]
  assign CAMLine_68_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_68_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_69_clock = clock;
  assign CAMLine_69_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_69_io_wi = io_waddr[69]; // @[cam.scala 86:31]
  assign CAMLine_69_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_69_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_70_clock = clock;
  assign CAMLine_70_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_70_io_wi = io_waddr[70]; // @[cam.scala 86:31]
  assign CAMLine_70_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_70_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_71_clock = clock;
  assign CAMLine_71_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_71_io_wi = io_waddr[71]; // @[cam.scala 86:31]
  assign CAMLine_71_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_71_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_72_clock = clock;
  assign CAMLine_72_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_72_io_wi = io_waddr[72]; // @[cam.scala 86:31]
  assign CAMLine_72_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_72_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_73_clock = clock;
  assign CAMLine_73_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_73_io_wi = io_waddr[73]; // @[cam.scala 86:31]
  assign CAMLine_73_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_73_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_74_clock = clock;
  assign CAMLine_74_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_74_io_wi = io_waddr[74]; // @[cam.scala 86:31]
  assign CAMLine_74_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_74_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_75_clock = clock;
  assign CAMLine_75_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_75_io_wi = io_waddr[75]; // @[cam.scala 86:31]
  assign CAMLine_75_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_75_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_76_clock = clock;
  assign CAMLine_76_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_76_io_wi = io_waddr[76]; // @[cam.scala 86:31]
  assign CAMLine_76_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_76_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_77_clock = clock;
  assign CAMLine_77_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_77_io_wi = io_waddr[77]; // @[cam.scala 86:31]
  assign CAMLine_77_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_77_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_78_clock = clock;
  assign CAMLine_78_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_78_io_wi = io_waddr[78]; // @[cam.scala 86:31]
  assign CAMLine_78_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_78_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_79_clock = clock;
  assign CAMLine_79_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_79_io_wi = io_waddr[79]; // @[cam.scala 86:31]
  assign CAMLine_79_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_79_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_80_clock = clock;
  assign CAMLine_80_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_80_io_wi = io_waddr[80]; // @[cam.scala 86:31]
  assign CAMLine_80_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_80_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_81_clock = clock;
  assign CAMLine_81_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_81_io_wi = io_waddr[81]; // @[cam.scala 86:31]
  assign CAMLine_81_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_81_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_82_clock = clock;
  assign CAMLine_82_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_82_io_wi = io_waddr[82]; // @[cam.scala 86:31]
  assign CAMLine_82_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_82_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_83_clock = clock;
  assign CAMLine_83_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_83_io_wi = io_waddr[83]; // @[cam.scala 86:31]
  assign CAMLine_83_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_83_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_84_clock = clock;
  assign CAMLine_84_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_84_io_wi = io_waddr[84]; // @[cam.scala 86:31]
  assign CAMLine_84_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_84_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_85_clock = clock;
  assign CAMLine_85_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_85_io_wi = io_waddr[85]; // @[cam.scala 86:31]
  assign CAMLine_85_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_85_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_86_clock = clock;
  assign CAMLine_86_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_86_io_wi = io_waddr[86]; // @[cam.scala 86:31]
  assign CAMLine_86_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_86_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_87_clock = clock;
  assign CAMLine_87_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_87_io_wi = io_waddr[87]; // @[cam.scala 86:31]
  assign CAMLine_87_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_87_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_88_clock = clock;
  assign CAMLine_88_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_88_io_wi = io_waddr[88]; // @[cam.scala 86:31]
  assign CAMLine_88_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_88_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_89_clock = clock;
  assign CAMLine_89_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_89_io_wi = io_waddr[89]; // @[cam.scala 86:31]
  assign CAMLine_89_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_89_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_90_clock = clock;
  assign CAMLine_90_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_90_io_wi = io_waddr[90]; // @[cam.scala 86:31]
  assign CAMLine_90_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_90_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_91_clock = clock;
  assign CAMLine_91_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_91_io_wi = io_waddr[91]; // @[cam.scala 86:31]
  assign CAMLine_91_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_91_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_92_clock = clock;
  assign CAMLine_92_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_92_io_wi = io_waddr[92]; // @[cam.scala 86:31]
  assign CAMLine_92_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_92_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_93_clock = clock;
  assign CAMLine_93_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_93_io_wi = io_waddr[93]; // @[cam.scala 86:31]
  assign CAMLine_93_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_93_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_94_clock = clock;
  assign CAMLine_94_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_94_io_wi = io_waddr[94]; // @[cam.scala 86:31]
  assign CAMLine_94_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_94_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_95_clock = clock;
  assign CAMLine_95_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_95_io_wi = io_waddr[95]; // @[cam.scala 86:31]
  assign CAMLine_95_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_95_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_96_clock = clock;
  assign CAMLine_96_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_96_io_wi = io_waddr[96]; // @[cam.scala 86:31]
  assign CAMLine_96_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_96_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_97_clock = clock;
  assign CAMLine_97_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_97_io_wi = io_waddr[97]; // @[cam.scala 86:31]
  assign CAMLine_97_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_97_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_98_clock = clock;
  assign CAMLine_98_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_98_io_wi = io_waddr[98]; // @[cam.scala 86:31]
  assign CAMLine_98_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_98_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_99_clock = clock;
  assign CAMLine_99_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_99_io_wi = io_waddr[99]; // @[cam.scala 86:31]
  assign CAMLine_99_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_99_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_100_clock = clock;
  assign CAMLine_100_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_100_io_wi = io_waddr[100]; // @[cam.scala 86:31]
  assign CAMLine_100_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_100_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_101_clock = clock;
  assign CAMLine_101_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_101_io_wi = io_waddr[101]; // @[cam.scala 86:31]
  assign CAMLine_101_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_101_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_102_clock = clock;
  assign CAMLine_102_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_102_io_wi = io_waddr[102]; // @[cam.scala 86:31]
  assign CAMLine_102_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_102_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_103_clock = clock;
  assign CAMLine_103_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_103_io_wi = io_waddr[103]; // @[cam.scala 86:31]
  assign CAMLine_103_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_103_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_104_clock = clock;
  assign CAMLine_104_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_104_io_wi = io_waddr[104]; // @[cam.scala 86:31]
  assign CAMLine_104_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_104_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_105_clock = clock;
  assign CAMLine_105_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_105_io_wi = io_waddr[105]; // @[cam.scala 86:31]
  assign CAMLine_105_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_105_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_106_clock = clock;
  assign CAMLine_106_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_106_io_wi = io_waddr[106]; // @[cam.scala 86:31]
  assign CAMLine_106_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_106_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_107_clock = clock;
  assign CAMLine_107_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_107_io_wi = io_waddr[107]; // @[cam.scala 86:31]
  assign CAMLine_107_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_107_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_108_clock = clock;
  assign CAMLine_108_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_108_io_wi = io_waddr[108]; // @[cam.scala 86:31]
  assign CAMLine_108_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_108_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_109_clock = clock;
  assign CAMLine_109_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_109_io_wi = io_waddr[109]; // @[cam.scala 86:31]
  assign CAMLine_109_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_109_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_110_clock = clock;
  assign CAMLine_110_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_110_io_wi = io_waddr[110]; // @[cam.scala 86:31]
  assign CAMLine_110_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_110_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_111_clock = clock;
  assign CAMLine_111_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_111_io_wi = io_waddr[111]; // @[cam.scala 86:31]
  assign CAMLine_111_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_111_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_112_clock = clock;
  assign CAMLine_112_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_112_io_wi = io_waddr[112]; // @[cam.scala 86:31]
  assign CAMLine_112_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_112_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_113_clock = clock;
  assign CAMLine_113_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_113_io_wi = io_waddr[113]; // @[cam.scala 86:31]
  assign CAMLine_113_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_113_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_114_clock = clock;
  assign CAMLine_114_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_114_io_wi = io_waddr[114]; // @[cam.scala 86:31]
  assign CAMLine_114_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_114_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_115_clock = clock;
  assign CAMLine_115_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_115_io_wi = io_waddr[115]; // @[cam.scala 86:31]
  assign CAMLine_115_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_115_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_116_clock = clock;
  assign CAMLine_116_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_116_io_wi = io_waddr[116]; // @[cam.scala 86:31]
  assign CAMLine_116_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_116_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_117_clock = clock;
  assign CAMLine_117_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_117_io_wi = io_waddr[117]; // @[cam.scala 86:31]
  assign CAMLine_117_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_117_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_118_clock = clock;
  assign CAMLine_118_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_118_io_wi = io_waddr[118]; // @[cam.scala 86:31]
  assign CAMLine_118_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_118_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_119_clock = clock;
  assign CAMLine_119_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_119_io_wi = io_waddr[119]; // @[cam.scala 86:31]
  assign CAMLine_119_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_119_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_120_clock = clock;
  assign CAMLine_120_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_120_io_wi = io_waddr[120]; // @[cam.scala 86:31]
  assign CAMLine_120_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_120_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_121_clock = clock;
  assign CAMLine_121_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_121_io_wi = io_waddr[121]; // @[cam.scala 86:31]
  assign CAMLine_121_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_121_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_122_clock = clock;
  assign CAMLine_122_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_122_io_wi = io_waddr[122]; // @[cam.scala 86:31]
  assign CAMLine_122_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_122_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_123_clock = clock;
  assign CAMLine_123_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_123_io_wi = io_waddr[123]; // @[cam.scala 86:31]
  assign CAMLine_123_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_123_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_124_clock = clock;
  assign CAMLine_124_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_124_io_wi = io_waddr[124]; // @[cam.scala 86:31]
  assign CAMLine_124_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_124_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_125_clock = clock;
  assign CAMLine_125_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_125_io_wi = io_waddr[125]; // @[cam.scala 86:31]
  assign CAMLine_125_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_125_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_126_clock = clock;
  assign CAMLine_126_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_126_io_wi = io_waddr[126]; // @[cam.scala 86:31]
  assign CAMLine_126_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_126_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_127_clock = clock;
  assign CAMLine_127_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_127_io_wi = io_waddr[127]; // @[cam.scala 86:31]
  assign CAMLine_127_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_127_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_128_clock = clock;
  assign CAMLine_128_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_128_io_wi = io_waddr[128]; // @[cam.scala 86:31]
  assign CAMLine_128_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_128_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_129_clock = clock;
  assign CAMLine_129_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_129_io_wi = io_waddr[129]; // @[cam.scala 86:31]
  assign CAMLine_129_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_129_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_130_clock = clock;
  assign CAMLine_130_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_130_io_wi = io_waddr[130]; // @[cam.scala 86:31]
  assign CAMLine_130_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_130_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_131_clock = clock;
  assign CAMLine_131_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_131_io_wi = io_waddr[131]; // @[cam.scala 86:31]
  assign CAMLine_131_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_131_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_132_clock = clock;
  assign CAMLine_132_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_132_io_wi = io_waddr[132]; // @[cam.scala 86:31]
  assign CAMLine_132_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_132_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_133_clock = clock;
  assign CAMLine_133_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_133_io_wi = io_waddr[133]; // @[cam.scala 86:31]
  assign CAMLine_133_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_133_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_134_clock = clock;
  assign CAMLine_134_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_134_io_wi = io_waddr[134]; // @[cam.scala 86:31]
  assign CAMLine_134_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_134_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_135_clock = clock;
  assign CAMLine_135_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_135_io_wi = io_waddr[135]; // @[cam.scala 86:31]
  assign CAMLine_135_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_135_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_136_clock = clock;
  assign CAMLine_136_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_136_io_wi = io_waddr[136]; // @[cam.scala 86:31]
  assign CAMLine_136_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_136_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_137_clock = clock;
  assign CAMLine_137_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_137_io_wi = io_waddr[137]; // @[cam.scala 86:31]
  assign CAMLine_137_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_137_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_138_clock = clock;
  assign CAMLine_138_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_138_io_wi = io_waddr[138]; // @[cam.scala 86:31]
  assign CAMLine_138_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_138_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_139_clock = clock;
  assign CAMLine_139_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_139_io_wi = io_waddr[139]; // @[cam.scala 86:31]
  assign CAMLine_139_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_139_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_140_clock = clock;
  assign CAMLine_140_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_140_io_wi = io_waddr[140]; // @[cam.scala 86:31]
  assign CAMLine_140_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_140_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_141_clock = clock;
  assign CAMLine_141_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_141_io_wi = io_waddr[141]; // @[cam.scala 86:31]
  assign CAMLine_141_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_141_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_142_clock = clock;
  assign CAMLine_142_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_142_io_wi = io_waddr[142]; // @[cam.scala 86:31]
  assign CAMLine_142_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_142_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_143_clock = clock;
  assign CAMLine_143_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_143_io_wi = io_waddr[143]; // @[cam.scala 86:31]
  assign CAMLine_143_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_143_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_144_clock = clock;
  assign CAMLine_144_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_144_io_wi = io_waddr[144]; // @[cam.scala 86:31]
  assign CAMLine_144_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_144_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_145_clock = clock;
  assign CAMLine_145_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_145_io_wi = io_waddr[145]; // @[cam.scala 86:31]
  assign CAMLine_145_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_145_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_146_clock = clock;
  assign CAMLine_146_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_146_io_wi = io_waddr[146]; // @[cam.scala 86:31]
  assign CAMLine_146_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_146_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_147_clock = clock;
  assign CAMLine_147_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_147_io_wi = io_waddr[147]; // @[cam.scala 86:31]
  assign CAMLine_147_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_147_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_148_clock = clock;
  assign CAMLine_148_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_148_io_wi = io_waddr[148]; // @[cam.scala 86:31]
  assign CAMLine_148_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_148_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_149_clock = clock;
  assign CAMLine_149_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_149_io_wi = io_waddr[149]; // @[cam.scala 86:31]
  assign CAMLine_149_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_149_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_150_clock = clock;
  assign CAMLine_150_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_150_io_wi = io_waddr[150]; // @[cam.scala 86:31]
  assign CAMLine_150_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_150_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_151_clock = clock;
  assign CAMLine_151_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_151_io_wi = io_waddr[151]; // @[cam.scala 86:31]
  assign CAMLine_151_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_151_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_152_clock = clock;
  assign CAMLine_152_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_152_io_wi = io_waddr[152]; // @[cam.scala 86:31]
  assign CAMLine_152_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_152_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_153_clock = clock;
  assign CAMLine_153_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_153_io_wi = io_waddr[153]; // @[cam.scala 86:31]
  assign CAMLine_153_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_153_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_154_clock = clock;
  assign CAMLine_154_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_154_io_wi = io_waddr[154]; // @[cam.scala 86:31]
  assign CAMLine_154_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_154_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_155_clock = clock;
  assign CAMLine_155_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_155_io_wi = io_waddr[155]; // @[cam.scala 86:31]
  assign CAMLine_155_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_155_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_156_clock = clock;
  assign CAMLine_156_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_156_io_wi = io_waddr[156]; // @[cam.scala 86:31]
  assign CAMLine_156_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_156_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_157_clock = clock;
  assign CAMLine_157_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_157_io_wi = io_waddr[157]; // @[cam.scala 86:31]
  assign CAMLine_157_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_157_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_158_clock = clock;
  assign CAMLine_158_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_158_io_wi = io_waddr[158]; // @[cam.scala 86:31]
  assign CAMLine_158_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_158_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_159_clock = clock;
  assign CAMLine_159_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_159_io_wi = io_waddr[159]; // @[cam.scala 86:31]
  assign CAMLine_159_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_159_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_160_clock = clock;
  assign CAMLine_160_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_160_io_wi = io_waddr[160]; // @[cam.scala 86:31]
  assign CAMLine_160_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_160_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_161_clock = clock;
  assign CAMLine_161_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_161_io_wi = io_waddr[161]; // @[cam.scala 86:31]
  assign CAMLine_161_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_161_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_162_clock = clock;
  assign CAMLine_162_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_162_io_wi = io_waddr[162]; // @[cam.scala 86:31]
  assign CAMLine_162_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_162_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_163_clock = clock;
  assign CAMLine_163_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_163_io_wi = io_waddr[163]; // @[cam.scala 86:31]
  assign CAMLine_163_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_163_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_164_clock = clock;
  assign CAMLine_164_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_164_io_wi = io_waddr[164]; // @[cam.scala 86:31]
  assign CAMLine_164_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_164_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_165_clock = clock;
  assign CAMLine_165_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_165_io_wi = io_waddr[165]; // @[cam.scala 86:31]
  assign CAMLine_165_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_165_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_166_clock = clock;
  assign CAMLine_166_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_166_io_wi = io_waddr[166]; // @[cam.scala 86:31]
  assign CAMLine_166_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_166_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_167_clock = clock;
  assign CAMLine_167_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_167_io_wi = io_waddr[167]; // @[cam.scala 86:31]
  assign CAMLine_167_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_167_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_168_clock = clock;
  assign CAMLine_168_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_168_io_wi = io_waddr[168]; // @[cam.scala 86:31]
  assign CAMLine_168_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_168_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_169_clock = clock;
  assign CAMLine_169_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_169_io_wi = io_waddr[169]; // @[cam.scala 86:31]
  assign CAMLine_169_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_169_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_170_clock = clock;
  assign CAMLine_170_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_170_io_wi = io_waddr[170]; // @[cam.scala 86:31]
  assign CAMLine_170_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_170_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_171_clock = clock;
  assign CAMLine_171_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_171_io_wi = io_waddr[171]; // @[cam.scala 86:31]
  assign CAMLine_171_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_171_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_172_clock = clock;
  assign CAMLine_172_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_172_io_wi = io_waddr[172]; // @[cam.scala 86:31]
  assign CAMLine_172_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_172_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_173_clock = clock;
  assign CAMLine_173_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_173_io_wi = io_waddr[173]; // @[cam.scala 86:31]
  assign CAMLine_173_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_173_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_174_clock = clock;
  assign CAMLine_174_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_174_io_wi = io_waddr[174]; // @[cam.scala 86:31]
  assign CAMLine_174_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_174_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_175_clock = clock;
  assign CAMLine_175_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_175_io_wi = io_waddr[175]; // @[cam.scala 86:31]
  assign CAMLine_175_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_175_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_176_clock = clock;
  assign CAMLine_176_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_176_io_wi = io_waddr[176]; // @[cam.scala 86:31]
  assign CAMLine_176_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_176_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_177_clock = clock;
  assign CAMLine_177_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_177_io_wi = io_waddr[177]; // @[cam.scala 86:31]
  assign CAMLine_177_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_177_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_178_clock = clock;
  assign CAMLine_178_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_178_io_wi = io_waddr[178]; // @[cam.scala 86:31]
  assign CAMLine_178_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_178_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_179_clock = clock;
  assign CAMLine_179_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_179_io_wi = io_waddr[179]; // @[cam.scala 86:31]
  assign CAMLine_179_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_179_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_180_clock = clock;
  assign CAMLine_180_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_180_io_wi = io_waddr[180]; // @[cam.scala 86:31]
  assign CAMLine_180_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_180_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_181_clock = clock;
  assign CAMLine_181_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_181_io_wi = io_waddr[181]; // @[cam.scala 86:31]
  assign CAMLine_181_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_181_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_182_clock = clock;
  assign CAMLine_182_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_182_io_wi = io_waddr[182]; // @[cam.scala 86:31]
  assign CAMLine_182_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_182_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_183_clock = clock;
  assign CAMLine_183_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_183_io_wi = io_waddr[183]; // @[cam.scala 86:31]
  assign CAMLine_183_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_183_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_184_clock = clock;
  assign CAMLine_184_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_184_io_wi = io_waddr[184]; // @[cam.scala 86:31]
  assign CAMLine_184_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_184_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_185_clock = clock;
  assign CAMLine_185_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_185_io_wi = io_waddr[185]; // @[cam.scala 86:31]
  assign CAMLine_185_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_185_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_186_clock = clock;
  assign CAMLine_186_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_186_io_wi = io_waddr[186]; // @[cam.scala 86:31]
  assign CAMLine_186_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_186_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_187_clock = clock;
  assign CAMLine_187_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_187_io_wi = io_waddr[187]; // @[cam.scala 86:31]
  assign CAMLine_187_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_187_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_188_clock = clock;
  assign CAMLine_188_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_188_io_wi = io_waddr[188]; // @[cam.scala 86:31]
  assign CAMLine_188_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_188_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_189_clock = clock;
  assign CAMLine_189_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_189_io_wi = io_waddr[189]; // @[cam.scala 86:31]
  assign CAMLine_189_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_189_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_190_clock = clock;
  assign CAMLine_190_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_190_io_wi = io_waddr[190]; // @[cam.scala 86:31]
  assign CAMLine_190_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_190_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_191_clock = clock;
  assign CAMLine_191_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_191_io_wi = io_waddr[191]; // @[cam.scala 86:31]
  assign CAMLine_191_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_191_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_192_clock = clock;
  assign CAMLine_192_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_192_io_wi = io_waddr[192]; // @[cam.scala 86:31]
  assign CAMLine_192_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_192_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_193_clock = clock;
  assign CAMLine_193_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_193_io_wi = io_waddr[193]; // @[cam.scala 86:31]
  assign CAMLine_193_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_193_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_194_clock = clock;
  assign CAMLine_194_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_194_io_wi = io_waddr[194]; // @[cam.scala 86:31]
  assign CAMLine_194_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_194_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_195_clock = clock;
  assign CAMLine_195_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_195_io_wi = io_waddr[195]; // @[cam.scala 86:31]
  assign CAMLine_195_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_195_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_196_clock = clock;
  assign CAMLine_196_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_196_io_wi = io_waddr[196]; // @[cam.scala 86:31]
  assign CAMLine_196_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_196_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_197_clock = clock;
  assign CAMLine_197_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_197_io_wi = io_waddr[197]; // @[cam.scala 86:31]
  assign CAMLine_197_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_197_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_198_clock = clock;
  assign CAMLine_198_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_198_io_wi = io_waddr[198]; // @[cam.scala 86:31]
  assign CAMLine_198_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_198_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_199_clock = clock;
  assign CAMLine_199_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_199_io_wi = io_waddr[199]; // @[cam.scala 86:31]
  assign CAMLine_199_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_199_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_200_clock = clock;
  assign CAMLine_200_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_200_io_wi = io_waddr[200]; // @[cam.scala 86:31]
  assign CAMLine_200_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_200_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_201_clock = clock;
  assign CAMLine_201_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_201_io_wi = io_waddr[201]; // @[cam.scala 86:31]
  assign CAMLine_201_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_201_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_202_clock = clock;
  assign CAMLine_202_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_202_io_wi = io_waddr[202]; // @[cam.scala 86:31]
  assign CAMLine_202_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_202_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_203_clock = clock;
  assign CAMLine_203_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_203_io_wi = io_waddr[203]; // @[cam.scala 86:31]
  assign CAMLine_203_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_203_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_204_clock = clock;
  assign CAMLine_204_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_204_io_wi = io_waddr[204]; // @[cam.scala 86:31]
  assign CAMLine_204_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_204_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_205_clock = clock;
  assign CAMLine_205_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_205_io_wi = io_waddr[205]; // @[cam.scala 86:31]
  assign CAMLine_205_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_205_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_206_clock = clock;
  assign CAMLine_206_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_206_io_wi = io_waddr[206]; // @[cam.scala 86:31]
  assign CAMLine_206_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_206_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_207_clock = clock;
  assign CAMLine_207_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_207_io_wi = io_waddr[207]; // @[cam.scala 86:31]
  assign CAMLine_207_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_207_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_208_clock = clock;
  assign CAMLine_208_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_208_io_wi = io_waddr[208]; // @[cam.scala 86:31]
  assign CAMLine_208_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_208_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_209_clock = clock;
  assign CAMLine_209_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_209_io_wi = io_waddr[209]; // @[cam.scala 86:31]
  assign CAMLine_209_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_209_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_210_clock = clock;
  assign CAMLine_210_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_210_io_wi = io_waddr[210]; // @[cam.scala 86:31]
  assign CAMLine_210_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_210_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_211_clock = clock;
  assign CAMLine_211_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_211_io_wi = io_waddr[211]; // @[cam.scala 86:31]
  assign CAMLine_211_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_211_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_212_clock = clock;
  assign CAMLine_212_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_212_io_wi = io_waddr[212]; // @[cam.scala 86:31]
  assign CAMLine_212_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_212_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_213_clock = clock;
  assign CAMLine_213_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_213_io_wi = io_waddr[213]; // @[cam.scala 86:31]
  assign CAMLine_213_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_213_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_214_clock = clock;
  assign CAMLine_214_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_214_io_wi = io_waddr[214]; // @[cam.scala 86:31]
  assign CAMLine_214_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_214_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_215_clock = clock;
  assign CAMLine_215_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_215_io_wi = io_waddr[215]; // @[cam.scala 86:31]
  assign CAMLine_215_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_215_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_216_clock = clock;
  assign CAMLine_216_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_216_io_wi = io_waddr[216]; // @[cam.scala 86:31]
  assign CAMLine_216_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_216_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_217_clock = clock;
  assign CAMLine_217_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_217_io_wi = io_waddr[217]; // @[cam.scala 86:31]
  assign CAMLine_217_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_217_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_218_clock = clock;
  assign CAMLine_218_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_218_io_wi = io_waddr[218]; // @[cam.scala 86:31]
  assign CAMLine_218_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_218_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_219_clock = clock;
  assign CAMLine_219_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_219_io_wi = io_waddr[219]; // @[cam.scala 86:31]
  assign CAMLine_219_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_219_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_220_clock = clock;
  assign CAMLine_220_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_220_io_wi = io_waddr[220]; // @[cam.scala 86:31]
  assign CAMLine_220_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_220_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_221_clock = clock;
  assign CAMLine_221_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_221_io_wi = io_waddr[221]; // @[cam.scala 86:31]
  assign CAMLine_221_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_221_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_222_clock = clock;
  assign CAMLine_222_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_222_io_wi = io_waddr[222]; // @[cam.scala 86:31]
  assign CAMLine_222_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_222_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_223_clock = clock;
  assign CAMLine_223_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_223_io_wi = io_waddr[223]; // @[cam.scala 86:31]
  assign CAMLine_223_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_223_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_224_clock = clock;
  assign CAMLine_224_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_224_io_wi = io_waddr[224]; // @[cam.scala 86:31]
  assign CAMLine_224_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_224_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_225_clock = clock;
  assign CAMLine_225_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_225_io_wi = io_waddr[225]; // @[cam.scala 86:31]
  assign CAMLine_225_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_225_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_226_clock = clock;
  assign CAMLine_226_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_226_io_wi = io_waddr[226]; // @[cam.scala 86:31]
  assign CAMLine_226_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_226_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_227_clock = clock;
  assign CAMLine_227_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_227_io_wi = io_waddr[227]; // @[cam.scala 86:31]
  assign CAMLine_227_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_227_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_228_clock = clock;
  assign CAMLine_228_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_228_io_wi = io_waddr[228]; // @[cam.scala 86:31]
  assign CAMLine_228_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_228_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_229_clock = clock;
  assign CAMLine_229_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_229_io_wi = io_waddr[229]; // @[cam.scala 86:31]
  assign CAMLine_229_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_229_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_230_clock = clock;
  assign CAMLine_230_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_230_io_wi = io_waddr[230]; // @[cam.scala 86:31]
  assign CAMLine_230_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_230_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_231_clock = clock;
  assign CAMLine_231_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_231_io_wi = io_waddr[231]; // @[cam.scala 86:31]
  assign CAMLine_231_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_231_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_232_clock = clock;
  assign CAMLine_232_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_232_io_wi = io_waddr[232]; // @[cam.scala 86:31]
  assign CAMLine_232_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_232_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_233_clock = clock;
  assign CAMLine_233_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_233_io_wi = io_waddr[233]; // @[cam.scala 86:31]
  assign CAMLine_233_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_233_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_234_clock = clock;
  assign CAMLine_234_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_234_io_wi = io_waddr[234]; // @[cam.scala 86:31]
  assign CAMLine_234_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_234_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_235_clock = clock;
  assign CAMLine_235_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_235_io_wi = io_waddr[235]; // @[cam.scala 86:31]
  assign CAMLine_235_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_235_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_236_clock = clock;
  assign CAMLine_236_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_236_io_wi = io_waddr[236]; // @[cam.scala 86:31]
  assign CAMLine_236_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_236_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_237_clock = clock;
  assign CAMLine_237_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_237_io_wi = io_waddr[237]; // @[cam.scala 86:31]
  assign CAMLine_237_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_237_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_238_clock = clock;
  assign CAMLine_238_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_238_io_wi = io_waddr[238]; // @[cam.scala 86:31]
  assign CAMLine_238_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_238_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_239_clock = clock;
  assign CAMLine_239_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_239_io_wi = io_waddr[239]; // @[cam.scala 86:31]
  assign CAMLine_239_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_239_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_240_clock = clock;
  assign CAMLine_240_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_240_io_wi = io_waddr[240]; // @[cam.scala 86:31]
  assign CAMLine_240_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_240_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_241_clock = clock;
  assign CAMLine_241_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_241_io_wi = io_waddr[241]; // @[cam.scala 86:31]
  assign CAMLine_241_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_241_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_242_clock = clock;
  assign CAMLine_242_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_242_io_wi = io_waddr[242]; // @[cam.scala 86:31]
  assign CAMLine_242_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_242_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_243_clock = clock;
  assign CAMLine_243_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_243_io_wi = io_waddr[243]; // @[cam.scala 86:31]
  assign CAMLine_243_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_243_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_244_clock = clock;
  assign CAMLine_244_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_244_io_wi = io_waddr[244]; // @[cam.scala 86:31]
  assign CAMLine_244_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_244_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_245_clock = clock;
  assign CAMLine_245_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_245_io_wi = io_waddr[245]; // @[cam.scala 86:31]
  assign CAMLine_245_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_245_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_246_clock = clock;
  assign CAMLine_246_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_246_io_wi = io_waddr[246]; // @[cam.scala 86:31]
  assign CAMLine_246_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_246_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_247_clock = clock;
  assign CAMLine_247_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_247_io_wi = io_waddr[247]; // @[cam.scala 86:31]
  assign CAMLine_247_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_247_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_248_clock = clock;
  assign CAMLine_248_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_248_io_wi = io_waddr[248]; // @[cam.scala 86:31]
  assign CAMLine_248_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_248_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_249_clock = clock;
  assign CAMLine_249_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_249_io_wi = io_waddr[249]; // @[cam.scala 86:31]
  assign CAMLine_249_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_249_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_250_clock = clock;
  assign CAMLine_250_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_250_io_wi = io_waddr[250]; // @[cam.scala 86:31]
  assign CAMLine_250_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_250_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_251_clock = clock;
  assign CAMLine_251_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_251_io_wi = io_waddr[251]; // @[cam.scala 86:31]
  assign CAMLine_251_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_251_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_252_clock = clock;
  assign CAMLine_252_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_252_io_wi = io_waddr[252]; // @[cam.scala 86:31]
  assign CAMLine_252_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_252_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_253_clock = clock;
  assign CAMLine_253_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_253_io_wi = io_waddr[253]; // @[cam.scala 86:31]
  assign CAMLine_253_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_253_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_254_clock = clock;
  assign CAMLine_254_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_254_io_wi = io_waddr[254]; // @[cam.scala 86:31]
  assign CAMLine_254_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_254_io_din = io_din; // @[cam.scala 88:21]
  assign CAMLine_255_clock = clock;
  assign CAMLine_255_io_we = io_we; // @[cam.scala 85:20]
  assign CAMLine_255_io_wi = io_waddr[255]; // @[cam.scala 86:31]
  assign CAMLine_255_io_key = io_key; // @[cam.scala 87:21]
  assign CAMLine_255_io_din = io_din; // @[cam.scala 88:21]
endmodule
